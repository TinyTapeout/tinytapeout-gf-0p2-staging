VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_MichaelBell_tinyQV
  CLASS BLOCK ;
  FOREIGN tt_um_MichaelBell_tinyQV ;
  ORIGIN 0.000 0.000 ;
  SIZE 1075.760 BY 736.960 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.780 3.620 177.380 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.380 3.620 330.980 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 482.980 3.620 484.580 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.580 3.620 638.180 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.180 3.620 791.780 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.780 3.620 945.380 733.340 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.480 3.620 174.080 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.080 3.620 327.680 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 479.680 3.620 481.280 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 633.280 3.620 634.880 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 786.880 3.620 788.480 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.480 3.620 942.080 733.340 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 331.090 735.960 331.390 736.960 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 338.370 735.960 338.670 736.960 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.810 735.960 324.110 736.960 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 316.530 735.960 316.830 736.960 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 309.250 735.960 309.550 736.960 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 301.970 735.960 302.270 736.960 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 294.690 735.960 294.990 736.960 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 287.410 735.960 287.710 736.960 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 280.130 735.960 280.430 736.960 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 272.850 735.960 273.150 736.960 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 265.570 735.960 265.870 736.960 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 258.290 735.960 258.590 736.960 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 251.010 735.960 251.310 736.960 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 243.730 735.960 244.030 736.960 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 236.450 735.960 236.750 736.960 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 229.170 735.960 229.470 736.960 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 221.890 735.960 222.190 736.960 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 214.610 735.960 214.910 736.960 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 207.330 735.960 207.630 736.960 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 83.570 735.960 83.870 736.960 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.069600 ;
    PORT
      LAYER Metal4 ;
        RECT 76.290 735.960 76.590 736.960 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 69.010 735.960 69.310 736.960 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 61.730 735.960 62.030 736.960 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 54.450 735.960 54.750 736.960 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.816000 ;
    ANTENNADIFFAREA 2.069600 ;
    PORT
      LAYER Metal4 ;
        RECT 47.170 735.960 47.470 736.960 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 39.890 735.960 40.190 736.960 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 32.610 735.960 32.910 736.960 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 141.810 735.960 142.110 736.960 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.219200 ;
    PORT
      LAYER Metal4 ;
        RECT 134.530 735.960 134.830 736.960 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.219200 ;
    PORT
      LAYER Metal4 ;
        RECT 127.250 735.960 127.550 736.960 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 119.970 735.960 120.270 736.960 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.879200 ;
    PORT
      LAYER Metal4 ;
        RECT 112.690 735.960 112.990 736.960 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.219200 ;
    PORT
      LAYER Metal4 ;
        RECT 105.410 735.960 105.710 736.960 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal4 ;
        RECT 98.130 735.960 98.430 736.960 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.389000 ;
    PORT
      LAYER Metal4 ;
        RECT 90.850 735.960 91.150 736.960 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.028900 ;
    PORT
      LAYER Metal4 ;
        RECT 200.050 735.960 200.350 736.960 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 192.770 735.960 193.070 736.960 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal4 ;
        RECT 185.490 735.960 185.790 736.960 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal4 ;
        RECT 178.210 735.960 178.510 736.960 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal4 ;
        RECT 170.930 735.960 171.230 736.960 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.121800 ;
    PORT
      LAYER Metal4 ;
        RECT 163.650 735.960 163.950 736.960 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.219200 ;
    PORT
      LAYER Metal4 ;
        RECT 156.370 735.960 156.670 736.960 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.879200 ;
    PORT
      LAYER Metal4 ;
        RECT 149.090 735.960 149.390 736.960 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 1073.390 733.470 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 1072.960 733.340 ;
      LAYER Metal2 ;
        RECT 1.820 0.090 1072.260 736.870 ;
      LAYER Metal3 ;
        RECT 1.770 0.140 1072.310 736.820 ;
      LAYER Metal4 ;
        RECT 8.540 735.660 32.310 735.960 ;
        RECT 33.210 735.660 39.590 735.960 ;
        RECT 40.490 735.660 46.870 735.960 ;
        RECT 47.770 735.660 54.150 735.960 ;
        RECT 55.050 735.660 61.430 735.960 ;
        RECT 62.330 735.660 68.710 735.960 ;
        RECT 69.610 735.660 75.990 735.960 ;
        RECT 76.890 735.660 83.270 735.960 ;
        RECT 84.170 735.660 90.550 735.960 ;
        RECT 91.450 735.660 97.830 735.960 ;
        RECT 98.730 735.660 105.110 735.960 ;
        RECT 106.010 735.660 112.390 735.960 ;
        RECT 113.290 735.660 119.670 735.960 ;
        RECT 120.570 735.660 126.950 735.960 ;
        RECT 127.850 735.660 134.230 735.960 ;
        RECT 135.130 735.660 141.510 735.960 ;
        RECT 142.410 735.660 148.790 735.960 ;
        RECT 149.690 735.660 156.070 735.960 ;
        RECT 156.970 735.660 163.350 735.960 ;
        RECT 164.250 735.660 170.630 735.960 ;
        RECT 171.530 735.660 177.910 735.960 ;
        RECT 178.810 735.660 185.190 735.960 ;
        RECT 186.090 735.660 192.470 735.960 ;
        RECT 193.370 735.660 199.750 735.960 ;
        RECT 200.650 735.660 207.030 735.960 ;
        RECT 207.930 735.660 214.310 735.960 ;
        RECT 215.210 735.660 221.590 735.960 ;
        RECT 222.490 735.660 228.870 735.960 ;
        RECT 229.770 735.660 236.150 735.960 ;
        RECT 237.050 735.660 243.430 735.960 ;
        RECT 244.330 735.660 250.710 735.960 ;
        RECT 251.610 735.660 257.990 735.960 ;
        RECT 258.890 735.660 265.270 735.960 ;
        RECT 266.170 735.660 272.550 735.960 ;
        RECT 273.450 735.660 279.830 735.960 ;
        RECT 280.730 735.660 287.110 735.960 ;
        RECT 288.010 735.660 294.390 735.960 ;
        RECT 295.290 735.660 301.670 735.960 ;
        RECT 302.570 735.660 308.950 735.960 ;
        RECT 309.850 735.660 316.230 735.960 ;
        RECT 317.130 735.660 323.510 735.960 ;
        RECT 324.410 735.660 330.790 735.960 ;
        RECT 331.690 735.660 338.070 735.960 ;
        RECT 338.970 735.660 1067.780 735.960 ;
        RECT 8.540 733.640 1067.780 735.660 ;
        RECT 8.540 3.320 18.580 733.640 ;
        RECT 20.780 3.320 21.880 733.640 ;
        RECT 24.080 3.320 172.180 733.640 ;
        RECT 174.380 3.320 175.480 733.640 ;
        RECT 177.680 3.320 325.780 733.640 ;
        RECT 327.980 3.320 329.080 733.640 ;
        RECT 331.280 3.320 479.380 733.640 ;
        RECT 481.580 3.320 482.680 733.640 ;
        RECT 484.880 3.320 632.980 733.640 ;
        RECT 635.180 3.320 636.280 733.640 ;
        RECT 638.480 3.320 786.580 733.640 ;
        RECT 788.780 3.320 789.880 733.640 ;
        RECT 792.080 3.320 940.180 733.640 ;
        RECT 942.380 3.320 943.480 733.640 ;
        RECT 945.680 3.320 1067.780 733.640 ;
        RECT 8.540 0.650 1067.780 3.320 ;
  END
END tt_um_MichaelBell_tinyQV
END LIBRARY


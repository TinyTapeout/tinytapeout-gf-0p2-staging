module tt_um_factory_test (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire clknet_0_clk;
 wire \cnt[0] ;
 wire \cnt[1] ;
 wire \cnt[2] ;
 wire \cnt[3] ;
 wire \cnt[4] ;
 wire \cnt[5] ;
 wire \cnt[6] ;
 wire \cnt[7] ;
 wire rst_n_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _035_ (.I(\cnt[0] ),
    .ZN(_000_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _036_ (.I(net2),
    .ZN(_008_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _037_ (.I(net18),
    .ZN(_009_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _038_ (.I(\cnt[5] ),
    .ZN(_010_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _039_ (.I(net7),
    .ZN(_011_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _040_ (.A1(_008_),
    .A2(_009_),
    .ZN(uio_oe[7]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _041_ (.A1(net10),
    .A2(net18),
    .ZN(_012_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _042_ (.A1(_000_),
    .A2(uio_oe[7]),
    .B1(_012_),
    .B2(_008_),
    .ZN(uo_out[0]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _043_ (.A1(net2),
    .A2(\cnt[1] ),
    .Z(uio_out[1]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _044_ (.A1(_008_),
    .A2(net11),
    .B(uio_out[1]),
    .ZN(_013_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _045_ (.A1(net18),
    .A2(net3),
    .ZN(_014_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _046_ (.A1(net18),
    .A2(_013_),
    .B(_014_),
    .ZN(uo_out[1]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _047_ (.A1(net2),
    .A2(\cnt[2] ),
    .Z(uio_out[2]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _048_ (.A1(_008_),
    .A2(net12),
    .B(uio_out[2]),
    .ZN(_015_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _049_ (.A1(net19),
    .A2(net4),
    .ZN(_016_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _050_ (.A1(net18),
    .A2(_015_),
    .B(_016_),
    .ZN(uo_out[2]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _051_ (.A1(net2),
    .A2(\cnt[3] ),
    .Z(uio_out[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _052_ (.A1(_008_),
    .A2(net13),
    .B(uio_out[3]),
    .ZN(_017_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _053_ (.A1(net19),
    .A2(net5),
    .ZN(_018_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _054_ (.A1(net18),
    .A2(_017_),
    .B(_018_),
    .ZN(uo_out[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _055_ (.A1(net2),
    .A2(\cnt[4] ),
    .Z(uio_out[4]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _056_ (.A1(_008_),
    .A2(net14),
    .B(uio_out[4]),
    .ZN(_019_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _057_ (.A1(net19),
    .A2(net6),
    .ZN(_020_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _058_ (.A1(net18),
    .A2(_019_),
    .B(_020_),
    .ZN(uo_out[4]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _059_ (.A1(_008_),
    .A2(net15),
    .ZN(_021_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _060_ (.A1(net2),
    .A2(\cnt[5] ),
    .Z(uio_out[5]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _061_ (.A1(_009_),
    .A2(uio_out[5]),
    .ZN(_022_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _062_ (.A1(_009_),
    .A2(_011_),
    .B1(_021_),
    .B2(_022_),
    .ZN(uo_out[5]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _063_ (.A1(net2),
    .A2(\cnt[6] ),
    .Z(uio_out[6]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _064_ (.A1(_008_),
    .A2(net16),
    .B(uio_out[6]),
    .ZN(_023_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _065_ (.A1(net19),
    .A2(net8),
    .ZN(_024_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _066_ (.A1(net18),
    .A2(_023_),
    .B(_024_),
    .ZN(uo_out[6]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _067_ (.A1(net2),
    .A2(\cnt[7] ),
    .Z(uio_out[7]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _068_ (.A1(_008_),
    .A2(net17),
    .B(uio_out[7]),
    .ZN(_025_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _069_ (.A1(net19),
    .A2(net9),
    .ZN(_026_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _070_ (.A1(net18),
    .A2(_025_),
    .B(_026_),
    .ZN(uo_out[7]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _071_ (.A1(_000_),
    .A2(_008_),
    .ZN(uio_out[0]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _072_ (.A1(\cnt[0] ),
    .A2(\cnt[1] ),
    .Z(_001_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _073_ (.A1(\cnt[0] ),
    .A2(\cnt[1] ),
    .A3(\cnt[2] ),
    .Z(_027_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _074_ (.A1(\cnt[0] ),
    .A2(\cnt[1] ),
    .B(\cnt[2] ),
    .ZN(_028_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _075_ (.A1(_027_),
    .A2(_028_),
    .ZN(_002_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _076_ (.A1(\cnt[3] ),
    .A2(_027_),
    .ZN(_029_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _077_ (.A1(\cnt[3] ),
    .A2(_027_),
    .Z(_003_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _078_ (.A1(\cnt[3] ),
    .A2(\cnt[4] ),
    .A3(_027_),
    .ZN(_030_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _079_ (.A1(\cnt[4] ),
    .A2(_029_),
    .ZN(_004_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _080_ (.A1(\cnt[3] ),
    .A2(\cnt[4] ),
    .A3(\cnt[5] ),
    .Z(_031_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _081_ (.A1(_027_),
    .A2(_031_),
    .Z(_032_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _082_ (.A1(_010_),
    .A2(_030_),
    .B(_032_),
    .ZN(_005_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _083_ (.A1(\cnt[6] ),
    .A2(_027_),
    .A3(_031_),
    .ZN(_033_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _084_ (.A1(\cnt[6] ),
    .A2(_032_),
    .Z(_006_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _085_ (.A1(\cnt[7] ),
    .A2(_033_),
    .ZN(_007_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _086_ (.D(_000_),
    .RN(rst_n_i),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\cnt[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _087_ (.D(_001_),
    .RN(rst_n_i),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\cnt[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _088_ (.D(_002_),
    .RN(rst_n_i),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\cnt[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _089_ (.D(_003_),
    .RN(rst_n_i),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\cnt[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _090_ (.D(_004_),
    .RN(rst_n_i),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\cnt[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _091_ (.D(_005_),
    .RN(rst_n_i),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\cnt[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _092_ (.D(_006_),
    .RN(rst_n_i),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\cnt[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _093_ (.D(_007_),
    .RN(rst_n_i),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\cnt[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _094_ (.D(net20),
    .RN(net18),
    .CLK(clknet_1_1__leaf_clk),
    .Q(rst_n_i),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _096_ (.I(uio_oe[7]),
    .Z(uio_oe[0]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _097_ (.I(uio_oe[7]),
    .Z(uio_oe[1]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _098_ (.I(uio_oe[7]),
    .Z(uio_oe[2]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _099_ (.I(uio_oe[7]),
    .Z(uio_oe[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _100_ (.I(uio_oe[7]),
    .Z(uio_oe[4]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _101_ (.I(uio_oe[7]),
    .Z(uio_oe[5]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _102_ (.I(uio_oe[7]),
    .Z(uio_oe[6]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_39 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_40 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_41 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_42 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_43 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_44 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_45 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_46 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_47 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_48 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_49 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_50 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_51 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_52 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_53 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_54 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_55 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_56 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_57 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_58 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_59 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_60 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_61 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_62 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_63 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_64 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_65 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_66 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_67 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_68 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_69 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_70 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_71 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_72 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_73 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_74 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_75 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_76 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_77 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_78 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_79 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_80 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_81 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_82 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_83 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_84 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_85 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_86 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_87 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_88 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_89 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_95 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_96 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_97 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_98 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_99 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_103 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_109 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_110 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_111 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_113 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_114 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_115 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_116 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_117 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_118 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_119 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_120 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_121 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_122 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_123 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_124 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_125 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_126 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_127 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_128 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_129 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_130 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_131 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_132 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_133 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_134 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_135 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_136 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_137 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_138 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_139 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_140 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_141 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_142 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_143 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_144 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_145 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_146 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_147 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_148 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_149 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_150 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_151 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_152 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_153 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_154 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_155 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_156 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_157 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_158 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_159 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_160 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_161 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_162 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_163 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_164 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_165 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_166 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_167 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_168 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_169 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_170 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_171 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_172 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_173 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_174 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_175 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_176 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_177 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_178 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_179 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_180 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_181 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_182 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_183 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_184 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_185 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_186 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_187 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_188 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_189 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_190 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_191 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_192 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_193 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_194 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_195 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_196 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_197 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_198 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_199 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_200 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_201 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_202 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_203 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_204 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_205 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_206 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_207 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_208 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_209 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_210 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_211 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_212 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_213 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_214 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_215 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_216 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_217 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_218 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_219 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_220 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_221 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_222 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_223 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_224 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_225 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_226 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_227 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_228 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_229 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_230 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_231 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_232 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_233 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_234 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_235 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_236 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_237 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_238 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_239 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_240 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_241 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_242 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_243 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_244 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_245 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_246 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_247 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_248 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_249 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_250 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_251 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_252 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_253 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_254 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_255 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_256 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_257 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_258 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_259 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_260 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_261 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_262 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_263 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_264 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_265 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_266 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_267 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_268 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_269 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_270 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_271 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_272 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_273 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_274 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_275 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_276 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_277 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_278 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_279 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_280 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_281 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_282 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_283 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_284 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_285 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_286 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_287 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_288 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_289 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_290 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_291 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_292 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_293 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_294 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_295 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_296 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_297 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_298 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_299 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_300 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_301 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_302 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_303 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_304 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_305 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_306 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_307 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_308 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_309 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_310 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_311 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_312 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_313 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_314 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_315 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_316 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_317 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_318 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_319 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_320 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_321 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_322 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_323 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_324 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_325 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_326 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_327 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_328 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_329 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_330 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_331 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_332 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_333 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_334 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_335 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_336 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_337 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_338 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_339 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_340 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_341 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_342 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_343 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_344 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_345 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_346 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_347 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_348 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_349 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_350 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_351 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_352 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_353 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_354 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_355 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_356 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_357 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_358 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_359 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_360 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_361 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_362 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_363 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_364 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_365 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_366 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_367 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_368 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_369 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_370 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_371 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_372 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_373 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_374 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_375 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_376 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_377 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_378 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_379 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_380 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_381 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_382 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_383 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_384 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_385 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_386 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_387 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_388 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_389 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_390 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_391 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_392 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_393 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_394 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_395 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_396 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_397 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_398 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_399 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_400 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_401 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_402 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_403 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_404 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_405 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_406 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_407 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_409 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_410 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_411 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_412 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_413 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_414 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_416 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_417 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_418 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_419 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_420 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_421 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_422 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_423 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_424 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_425 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(rst_n),
    .Z(net1),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 input2 (.I(ui_in[0]),
    .Z(net2),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(ui_in[1]),
    .Z(net3),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(ui_in[2]),
    .Z(net4),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(ui_in[3]),
    .Z(net5),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(ui_in[4]),
    .Z(net6),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(ui_in[5]),
    .Z(net7),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(ui_in[6]),
    .Z(net8),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(ui_in[7]),
    .Z(net9),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(uio_in[0]),
    .Z(net10),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(uio_in[1]),
    .Z(net11),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(uio_in[2]),
    .Z(net12),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(uio_in[3]),
    .Z(net13),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(uio_in[4]),
    .Z(net14),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(uio_in[5]),
    .Z(net15),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(uio_in[6]),
    .Z(net16),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(uio_in[7]),
    .Z(net17),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 fanout18 (.I(net1),
    .Z(net18),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout19 (.I(net1),
    .Z(net19),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tieh _094__20 (.Z(net20),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkload0 (.I(clknet_1_1__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_596 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_368 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_372 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_374 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_385 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_407 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_415 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_440 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_341 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_435 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_467 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_483 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_487 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_447 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_477 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_290 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_294 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_441 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_458 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_71 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_86 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_102 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_303 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_336 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_494 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_496 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_503 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_519 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_535 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_574 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_50 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_54 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_80 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_82 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_188 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_332 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_484 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_516 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_576 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_600 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_36 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_70 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_316 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_320 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_322 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_434 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_596 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
endmodule

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_MichaelBell_tinyQV
  CLASS BLOCK ;
  FOREIGN tt_um_MichaelBell_tinyQV ;
  ORIGIN 0.000 0.000 ;
  SIZE 1075.760 BY 736.960 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.780 3.620 177.380 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.380 3.620 330.980 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 482.980 3.620 484.580 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.580 3.620 638.180 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.180 3.620 791.780 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.780 3.620 945.380 733.340 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.480 3.620 174.080 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.080 3.620 327.680 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 479.680 3.620 481.280 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 633.280 3.620 634.880 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 786.880 3.620 788.480 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.480 3.620 942.080 733.340 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 331.090 735.960 331.390 736.960 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 338.370 735.960 338.670 736.960 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.810 735.960 324.110 736.960 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 316.530 735.960 316.830 736.960 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 309.250 735.960 309.550 736.960 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 301.970 735.960 302.270 736.960 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 294.690 735.960 294.990 736.960 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 287.410 735.960 287.710 736.960 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 280.130 735.960 280.430 736.960 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 272.850 735.960 273.150 736.960 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 265.570 735.960 265.870 736.960 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 258.290 735.960 258.590 736.960 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 251.010 735.960 251.310 736.960 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 243.730 735.960 244.030 736.960 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 236.450 735.960 236.750 736.960 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    PORT
      LAYER Metal4 ;
        RECT 229.170 735.960 229.470 736.960 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 221.890 735.960 222.190 736.960 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 214.610 735.960 214.910 736.960 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 207.330 735.960 207.630 736.960 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 83.570 735.960 83.870 736.960 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.071900 ;
    PORT
      LAYER Metal4 ;
        RECT 76.290 735.960 76.590 736.960 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 69.010 735.960 69.310 736.960 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 61.730 735.960 62.030 736.960 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 54.450 735.960 54.750 736.960 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 2.069600 ;
    PORT
      LAYER Metal4 ;
        RECT 47.170 735.960 47.470 736.960 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 39.890 735.960 40.190 736.960 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 32.610 735.960 32.910 736.960 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 141.810 735.960 142.110 736.960 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 134.530 735.960 134.830 736.960 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 127.250 735.960 127.550 736.960 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 119.970 735.960 120.270 736.960 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.932000 ;
    PORT
      LAYER Metal4 ;
        RECT 112.690 735.960 112.990 736.960 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 105.410 735.960 105.710 736.960 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 98.130 735.960 98.430 736.960 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.389000 ;
    PORT
      LAYER Metal4 ;
        RECT 90.850 735.960 91.150 736.960 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 200.050 735.960 200.350 736.960 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 192.770 735.960 193.070 736.960 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal4 ;
        RECT 185.490 735.960 185.790 736.960 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal4 ;
        RECT 178.210 735.960 178.510 736.960 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal4 ;
        RECT 170.930 735.960 171.230 736.960 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal4 ;
        RECT 163.650 735.960 163.950 736.960 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 156.370 735.960 156.670 736.960 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 149.090 735.960 149.390 736.960 ;
    END
  END uo_out[7]
  OBS
      LAYER Pwell ;
        RECT 2.930 731.280 1073.390 733.470 ;
      LAYER Nwell ;
        RECT 2.930 726.960 1073.390 731.280 ;
      LAYER Pwell ;
        RECT 2.930 723.440 1073.390 726.960 ;
      LAYER Nwell ;
        RECT 2.930 719.120 1073.390 723.440 ;
      LAYER Pwell ;
        RECT 2.930 715.600 1073.390 719.120 ;
      LAYER Nwell ;
        RECT 2.930 711.280 1073.390 715.600 ;
      LAYER Pwell ;
        RECT 2.930 707.760 1073.390 711.280 ;
      LAYER Nwell ;
        RECT 2.930 703.440 1073.390 707.760 ;
      LAYER Pwell ;
        RECT 2.930 699.920 1073.390 703.440 ;
      LAYER Nwell ;
        RECT 2.930 695.600 1073.390 699.920 ;
      LAYER Pwell ;
        RECT 2.930 692.080 1073.390 695.600 ;
      LAYER Nwell ;
        RECT 2.930 687.760 1073.390 692.080 ;
      LAYER Pwell ;
        RECT 2.930 684.240 1073.390 687.760 ;
      LAYER Nwell ;
        RECT 2.930 679.920 1073.390 684.240 ;
      LAYER Pwell ;
        RECT 2.930 676.400 1073.390 679.920 ;
      LAYER Nwell ;
        RECT 2.930 672.080 1073.390 676.400 ;
      LAYER Pwell ;
        RECT 2.930 668.560 1073.390 672.080 ;
      LAYER Nwell ;
        RECT 2.930 664.240 1073.390 668.560 ;
      LAYER Pwell ;
        RECT 2.930 660.720 1073.390 664.240 ;
      LAYER Nwell ;
        RECT 2.930 656.400 1073.390 660.720 ;
      LAYER Pwell ;
        RECT 2.930 652.880 1073.390 656.400 ;
      LAYER Nwell ;
        RECT 2.930 648.560 1073.390 652.880 ;
      LAYER Pwell ;
        RECT 2.930 645.040 1073.390 648.560 ;
      LAYER Nwell ;
        RECT 2.930 640.720 1073.390 645.040 ;
      LAYER Pwell ;
        RECT 2.930 637.200 1073.390 640.720 ;
      LAYER Nwell ;
        RECT 2.930 632.880 1073.390 637.200 ;
      LAYER Pwell ;
        RECT 2.930 629.360 1073.390 632.880 ;
      LAYER Nwell ;
        RECT 2.930 625.040 1073.390 629.360 ;
      LAYER Pwell ;
        RECT 2.930 621.520 1073.390 625.040 ;
      LAYER Nwell ;
        RECT 2.930 617.200 1073.390 621.520 ;
      LAYER Pwell ;
        RECT 2.930 613.680 1073.390 617.200 ;
      LAYER Nwell ;
        RECT 2.930 609.360 1073.390 613.680 ;
      LAYER Pwell ;
        RECT 2.930 605.840 1073.390 609.360 ;
      LAYER Nwell ;
        RECT 2.930 601.520 1073.390 605.840 ;
      LAYER Pwell ;
        RECT 2.930 598.000 1073.390 601.520 ;
      LAYER Nwell ;
        RECT 2.930 593.680 1073.390 598.000 ;
      LAYER Pwell ;
        RECT 2.930 590.160 1073.390 593.680 ;
      LAYER Nwell ;
        RECT 2.930 585.840 1073.390 590.160 ;
      LAYER Pwell ;
        RECT 2.930 582.320 1073.390 585.840 ;
      LAYER Nwell ;
        RECT 2.930 578.000 1073.390 582.320 ;
      LAYER Pwell ;
        RECT 2.930 574.480 1073.390 578.000 ;
      LAYER Nwell ;
        RECT 2.930 570.160 1073.390 574.480 ;
      LAYER Pwell ;
        RECT 2.930 566.640 1073.390 570.160 ;
      LAYER Nwell ;
        RECT 2.930 562.320 1073.390 566.640 ;
      LAYER Pwell ;
        RECT 2.930 558.800 1073.390 562.320 ;
      LAYER Nwell ;
        RECT 2.930 554.480 1073.390 558.800 ;
      LAYER Pwell ;
        RECT 2.930 550.960 1073.390 554.480 ;
      LAYER Nwell ;
        RECT 2.930 546.640 1073.390 550.960 ;
      LAYER Pwell ;
        RECT 2.930 543.120 1073.390 546.640 ;
      LAYER Nwell ;
        RECT 2.930 538.800 1073.390 543.120 ;
      LAYER Pwell ;
        RECT 2.930 535.280 1073.390 538.800 ;
      LAYER Nwell ;
        RECT 2.930 530.960 1073.390 535.280 ;
      LAYER Pwell ;
        RECT 2.930 527.440 1073.390 530.960 ;
      LAYER Nwell ;
        RECT 2.930 523.120 1073.390 527.440 ;
      LAYER Pwell ;
        RECT 2.930 519.600 1073.390 523.120 ;
      LAYER Nwell ;
        RECT 2.930 515.280 1073.390 519.600 ;
      LAYER Pwell ;
        RECT 2.930 511.760 1073.390 515.280 ;
      LAYER Nwell ;
        RECT 2.930 507.440 1073.390 511.760 ;
      LAYER Pwell ;
        RECT 2.930 503.920 1073.390 507.440 ;
      LAYER Nwell ;
        RECT 2.930 499.600 1073.390 503.920 ;
      LAYER Pwell ;
        RECT 2.930 496.080 1073.390 499.600 ;
      LAYER Nwell ;
        RECT 2.930 491.760 1073.390 496.080 ;
      LAYER Pwell ;
        RECT 2.930 488.240 1073.390 491.760 ;
      LAYER Nwell ;
        RECT 2.930 483.920 1073.390 488.240 ;
      LAYER Pwell ;
        RECT 2.930 480.400 1073.390 483.920 ;
      LAYER Nwell ;
        RECT 2.930 476.080 1073.390 480.400 ;
      LAYER Pwell ;
        RECT 2.930 472.560 1073.390 476.080 ;
      LAYER Nwell ;
        RECT 2.930 468.240 1073.390 472.560 ;
      LAYER Pwell ;
        RECT 2.930 464.720 1073.390 468.240 ;
      LAYER Nwell ;
        RECT 2.930 460.400 1073.390 464.720 ;
      LAYER Pwell ;
        RECT 2.930 456.880 1073.390 460.400 ;
      LAYER Nwell ;
        RECT 2.930 452.560 1073.390 456.880 ;
      LAYER Pwell ;
        RECT 2.930 449.040 1073.390 452.560 ;
      LAYER Nwell ;
        RECT 2.930 444.720 1073.390 449.040 ;
      LAYER Pwell ;
        RECT 2.930 441.200 1073.390 444.720 ;
      LAYER Nwell ;
        RECT 2.930 436.880 1073.390 441.200 ;
      LAYER Pwell ;
        RECT 2.930 433.360 1073.390 436.880 ;
      LAYER Nwell ;
        RECT 2.930 429.040 1073.390 433.360 ;
      LAYER Pwell ;
        RECT 2.930 425.520 1073.390 429.040 ;
      LAYER Nwell ;
        RECT 2.930 421.200 1073.390 425.520 ;
      LAYER Pwell ;
        RECT 2.930 417.680 1073.390 421.200 ;
      LAYER Nwell ;
        RECT 2.930 413.360 1073.390 417.680 ;
      LAYER Pwell ;
        RECT 2.930 409.840 1073.390 413.360 ;
      LAYER Nwell ;
        RECT 2.930 405.520 1073.390 409.840 ;
      LAYER Pwell ;
        RECT 2.930 402.000 1073.390 405.520 ;
      LAYER Nwell ;
        RECT 2.930 397.680 1073.390 402.000 ;
      LAYER Pwell ;
        RECT 2.930 394.160 1073.390 397.680 ;
      LAYER Nwell ;
        RECT 2.930 389.840 1073.390 394.160 ;
      LAYER Pwell ;
        RECT 2.930 386.320 1073.390 389.840 ;
      LAYER Nwell ;
        RECT 2.930 382.000 1073.390 386.320 ;
      LAYER Pwell ;
        RECT 2.930 378.480 1073.390 382.000 ;
      LAYER Nwell ;
        RECT 2.930 374.160 1073.390 378.480 ;
      LAYER Pwell ;
        RECT 2.930 370.640 1073.390 374.160 ;
      LAYER Nwell ;
        RECT 2.930 366.320 1073.390 370.640 ;
      LAYER Pwell ;
        RECT 2.930 362.800 1073.390 366.320 ;
      LAYER Nwell ;
        RECT 2.930 358.480 1073.390 362.800 ;
      LAYER Pwell ;
        RECT 2.930 354.960 1073.390 358.480 ;
      LAYER Nwell ;
        RECT 2.930 350.640 1073.390 354.960 ;
      LAYER Pwell ;
        RECT 2.930 347.120 1073.390 350.640 ;
      LAYER Nwell ;
        RECT 2.930 342.800 1073.390 347.120 ;
      LAYER Pwell ;
        RECT 2.930 339.280 1073.390 342.800 ;
      LAYER Nwell ;
        RECT 2.930 334.960 1073.390 339.280 ;
      LAYER Pwell ;
        RECT 2.930 331.440 1073.390 334.960 ;
      LAYER Nwell ;
        RECT 2.930 327.120 1073.390 331.440 ;
      LAYER Pwell ;
        RECT 2.930 323.600 1073.390 327.120 ;
      LAYER Nwell ;
        RECT 2.930 319.280 1073.390 323.600 ;
      LAYER Pwell ;
        RECT 2.930 315.760 1073.390 319.280 ;
      LAYER Nwell ;
        RECT 2.930 311.440 1073.390 315.760 ;
      LAYER Pwell ;
        RECT 2.930 307.920 1073.390 311.440 ;
      LAYER Nwell ;
        RECT 2.930 303.600 1073.390 307.920 ;
      LAYER Pwell ;
        RECT 2.930 300.080 1073.390 303.600 ;
      LAYER Nwell ;
        RECT 2.930 295.760 1073.390 300.080 ;
      LAYER Pwell ;
        RECT 2.930 292.240 1073.390 295.760 ;
      LAYER Nwell ;
        RECT 2.930 287.920 1073.390 292.240 ;
      LAYER Pwell ;
        RECT 2.930 284.400 1073.390 287.920 ;
      LAYER Nwell ;
        RECT 2.930 280.080 1073.390 284.400 ;
      LAYER Pwell ;
        RECT 2.930 276.560 1073.390 280.080 ;
      LAYER Nwell ;
        RECT 2.930 272.240 1073.390 276.560 ;
      LAYER Pwell ;
        RECT 2.930 268.720 1073.390 272.240 ;
      LAYER Nwell ;
        RECT 2.930 264.400 1073.390 268.720 ;
      LAYER Pwell ;
        RECT 2.930 260.880 1073.390 264.400 ;
      LAYER Nwell ;
        RECT 2.930 256.560 1073.390 260.880 ;
      LAYER Pwell ;
        RECT 2.930 253.040 1073.390 256.560 ;
      LAYER Nwell ;
        RECT 2.930 248.720 1073.390 253.040 ;
      LAYER Pwell ;
        RECT 2.930 245.200 1073.390 248.720 ;
      LAYER Nwell ;
        RECT 2.930 240.880 1073.390 245.200 ;
      LAYER Pwell ;
        RECT 2.930 237.360 1073.390 240.880 ;
      LAYER Nwell ;
        RECT 2.930 233.040 1073.390 237.360 ;
      LAYER Pwell ;
        RECT 2.930 229.520 1073.390 233.040 ;
      LAYER Nwell ;
        RECT 2.930 225.200 1073.390 229.520 ;
      LAYER Pwell ;
        RECT 2.930 221.680 1073.390 225.200 ;
      LAYER Nwell ;
        RECT 2.930 217.360 1073.390 221.680 ;
      LAYER Pwell ;
        RECT 2.930 213.840 1073.390 217.360 ;
      LAYER Nwell ;
        RECT 2.930 209.520 1073.390 213.840 ;
      LAYER Pwell ;
        RECT 2.930 206.000 1073.390 209.520 ;
      LAYER Nwell ;
        RECT 2.930 201.680 1073.390 206.000 ;
      LAYER Pwell ;
        RECT 2.930 198.160 1073.390 201.680 ;
      LAYER Nwell ;
        RECT 2.930 193.840 1073.390 198.160 ;
      LAYER Pwell ;
        RECT 2.930 190.320 1073.390 193.840 ;
      LAYER Nwell ;
        RECT 2.930 186.000 1073.390 190.320 ;
      LAYER Pwell ;
        RECT 2.930 182.480 1073.390 186.000 ;
      LAYER Nwell ;
        RECT 2.930 178.160 1073.390 182.480 ;
      LAYER Pwell ;
        RECT 2.930 174.640 1073.390 178.160 ;
      LAYER Nwell ;
        RECT 2.930 170.320 1073.390 174.640 ;
      LAYER Pwell ;
        RECT 2.930 166.800 1073.390 170.320 ;
      LAYER Nwell ;
        RECT 2.930 162.480 1073.390 166.800 ;
      LAYER Pwell ;
        RECT 2.930 158.960 1073.390 162.480 ;
      LAYER Nwell ;
        RECT 2.930 154.640 1073.390 158.960 ;
      LAYER Pwell ;
        RECT 2.930 151.120 1073.390 154.640 ;
      LAYER Nwell ;
        RECT 2.930 146.800 1073.390 151.120 ;
      LAYER Pwell ;
        RECT 2.930 143.280 1073.390 146.800 ;
      LAYER Nwell ;
        RECT 2.930 138.960 1073.390 143.280 ;
      LAYER Pwell ;
        RECT 2.930 135.440 1073.390 138.960 ;
      LAYER Nwell ;
        RECT 2.930 131.120 1073.390 135.440 ;
      LAYER Pwell ;
        RECT 2.930 127.600 1073.390 131.120 ;
      LAYER Nwell ;
        RECT 2.930 123.280 1073.390 127.600 ;
      LAYER Pwell ;
        RECT 2.930 119.760 1073.390 123.280 ;
      LAYER Nwell ;
        RECT 2.930 115.440 1073.390 119.760 ;
      LAYER Pwell ;
        RECT 2.930 111.920 1073.390 115.440 ;
      LAYER Nwell ;
        RECT 2.930 107.600 1073.390 111.920 ;
      LAYER Pwell ;
        RECT 2.930 104.080 1073.390 107.600 ;
      LAYER Nwell ;
        RECT 2.930 99.760 1073.390 104.080 ;
      LAYER Pwell ;
        RECT 2.930 96.240 1073.390 99.760 ;
      LAYER Nwell ;
        RECT 2.930 91.920 1073.390 96.240 ;
      LAYER Pwell ;
        RECT 2.930 88.400 1073.390 91.920 ;
      LAYER Nwell ;
        RECT 2.930 84.080 1073.390 88.400 ;
      LAYER Pwell ;
        RECT 2.930 80.560 1073.390 84.080 ;
      LAYER Nwell ;
        RECT 2.930 76.240 1073.390 80.560 ;
      LAYER Pwell ;
        RECT 2.930 72.720 1073.390 76.240 ;
      LAYER Nwell ;
        RECT 2.930 68.400 1073.390 72.720 ;
      LAYER Pwell ;
        RECT 2.930 64.880 1073.390 68.400 ;
      LAYER Nwell ;
        RECT 2.930 60.560 1073.390 64.880 ;
      LAYER Pwell ;
        RECT 2.930 57.040 1073.390 60.560 ;
      LAYER Nwell ;
        RECT 2.930 52.720 1073.390 57.040 ;
      LAYER Pwell ;
        RECT 2.930 49.200 1073.390 52.720 ;
      LAYER Nwell ;
        RECT 2.930 44.880 1073.390 49.200 ;
      LAYER Pwell ;
        RECT 2.930 41.360 1073.390 44.880 ;
      LAYER Nwell ;
        RECT 2.930 37.040 1073.390 41.360 ;
      LAYER Pwell ;
        RECT 2.930 33.520 1073.390 37.040 ;
      LAYER Nwell ;
        RECT 2.930 29.200 1073.390 33.520 ;
      LAYER Pwell ;
        RECT 2.930 25.680 1073.390 29.200 ;
      LAYER Nwell ;
        RECT 2.930 21.360 1073.390 25.680 ;
      LAYER Pwell ;
        RECT 2.930 17.840 1073.390 21.360 ;
      LAYER Nwell ;
        RECT 2.930 13.520 1073.390 17.840 ;
      LAYER Pwell ;
        RECT 2.930 10.000 1073.390 13.520 ;
      LAYER Nwell ;
        RECT 2.930 5.680 1073.390 10.000 ;
      LAYER Pwell ;
        RECT 2.930 3.490 1073.390 5.680 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 1072.960 733.340 ;
      LAYER Metal2 ;
        RECT 3.500 0.090 1071.700 733.230 ;
      LAYER Metal3 ;
        RECT 3.450 0.140 1071.750 733.180 ;
      LAYER Metal4 ;
        RECT 16.380 735.660 32.310 735.960 ;
        RECT 33.210 735.660 39.590 735.960 ;
        RECT 40.490 735.660 46.870 735.960 ;
        RECT 47.770 735.660 54.150 735.960 ;
        RECT 55.050 735.660 61.430 735.960 ;
        RECT 62.330 735.660 68.710 735.960 ;
        RECT 69.610 735.660 75.990 735.960 ;
        RECT 76.890 735.660 83.270 735.960 ;
        RECT 84.170 735.660 90.550 735.960 ;
        RECT 91.450 735.660 97.830 735.960 ;
        RECT 98.730 735.660 105.110 735.960 ;
        RECT 106.010 735.660 112.390 735.960 ;
        RECT 113.290 735.660 119.670 735.960 ;
        RECT 120.570 735.660 126.950 735.960 ;
        RECT 127.850 735.660 134.230 735.960 ;
        RECT 135.130 735.660 141.510 735.960 ;
        RECT 142.410 735.660 148.790 735.960 ;
        RECT 149.690 735.660 156.070 735.960 ;
        RECT 156.970 735.660 163.350 735.960 ;
        RECT 164.250 735.660 170.630 735.960 ;
        RECT 171.530 735.660 177.910 735.960 ;
        RECT 178.810 735.660 185.190 735.960 ;
        RECT 186.090 735.660 192.470 735.960 ;
        RECT 193.370 735.660 199.750 735.960 ;
        RECT 200.650 735.660 207.030 735.960 ;
        RECT 207.930 735.660 214.310 735.960 ;
        RECT 215.210 735.660 221.590 735.960 ;
        RECT 222.490 735.660 228.870 735.960 ;
        RECT 229.770 735.660 236.150 735.960 ;
        RECT 237.050 735.660 243.430 735.960 ;
        RECT 244.330 735.660 250.710 735.960 ;
        RECT 251.610 735.660 257.990 735.960 ;
        RECT 258.890 735.660 265.270 735.960 ;
        RECT 266.170 735.660 272.550 735.960 ;
        RECT 273.450 735.660 279.830 735.960 ;
        RECT 280.730 735.660 287.110 735.960 ;
        RECT 288.010 735.660 294.390 735.960 ;
        RECT 295.290 735.660 301.670 735.960 ;
        RECT 302.570 735.660 308.950 735.960 ;
        RECT 309.850 735.660 316.230 735.960 ;
        RECT 317.130 735.660 323.510 735.960 ;
        RECT 324.410 735.660 330.790 735.960 ;
        RECT 331.690 735.660 338.070 735.960 ;
        RECT 338.970 735.660 1065.540 735.960 ;
        RECT 16.380 733.640 1065.540 735.660 ;
        RECT 16.380 3.320 18.580 733.640 ;
        RECT 20.780 3.320 21.880 733.640 ;
        RECT 24.080 3.320 172.180 733.640 ;
        RECT 174.380 3.320 175.480 733.640 ;
        RECT 177.680 3.320 325.780 733.640 ;
        RECT 327.980 3.320 329.080 733.640 ;
        RECT 331.280 3.320 479.380 733.640 ;
        RECT 481.580 3.320 482.680 733.640 ;
        RECT 484.880 3.320 632.980 733.640 ;
        RECT 635.180 3.320 636.280 733.640 ;
        RECT 638.480 3.320 786.580 733.640 ;
        RECT 788.780 3.320 789.880 733.640 ;
        RECT 792.080 3.320 940.180 733.640 ;
        RECT 942.380 3.320 943.480 733.640 ;
        RECT 945.680 3.320 1065.540 733.640 ;
        RECT 16.380 0.650 1065.540 3.320 ;
  END
END tt_um_MichaelBell_tinyQV
END LIBRARY


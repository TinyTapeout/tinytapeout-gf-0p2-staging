module tt_um_calonso88_spi_i2c_reg_bank (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire i2c_sda_oe;
 wire spi_miso;
 wire \sunrise_digital_top_i.cpha_sync ;
 wire \sunrise_digital_top_i.cpol_sync ;
 wire \sunrise_digital_top_i.protrocol_sel_sync ;
 wire \sunrise_digital_top_i.rw_regs[0] ;
 wire \sunrise_digital_top_i.rw_regs[10] ;
 wire \sunrise_digital_top_i.rw_regs[11] ;
 wire \sunrise_digital_top_i.rw_regs[12] ;
 wire \sunrise_digital_top_i.rw_regs[13] ;
 wire \sunrise_digital_top_i.rw_regs[14] ;
 wire \sunrise_digital_top_i.rw_regs[15] ;
 wire \sunrise_digital_top_i.rw_regs[16] ;
 wire \sunrise_digital_top_i.rw_regs[17] ;
 wire \sunrise_digital_top_i.rw_regs[18] ;
 wire \sunrise_digital_top_i.rw_regs[19] ;
 wire \sunrise_digital_top_i.rw_regs[1] ;
 wire \sunrise_digital_top_i.rw_regs[20] ;
 wire \sunrise_digital_top_i.rw_regs[21] ;
 wire \sunrise_digital_top_i.rw_regs[22] ;
 wire \sunrise_digital_top_i.rw_regs[23] ;
 wire \sunrise_digital_top_i.rw_regs[24] ;
 wire \sunrise_digital_top_i.rw_regs[25] ;
 wire \sunrise_digital_top_i.rw_regs[26] ;
 wire \sunrise_digital_top_i.rw_regs[27] ;
 wire \sunrise_digital_top_i.rw_regs[28] ;
 wire \sunrise_digital_top_i.rw_regs[29] ;
 wire \sunrise_digital_top_i.rw_regs[2] ;
 wire \sunrise_digital_top_i.rw_regs[30] ;
 wire \sunrise_digital_top_i.rw_regs[31] ;
 wire \sunrise_digital_top_i.rw_regs[32] ;
 wire \sunrise_digital_top_i.rw_regs[33] ;
 wire \sunrise_digital_top_i.rw_regs[34] ;
 wire \sunrise_digital_top_i.rw_regs[35] ;
 wire \sunrise_digital_top_i.rw_regs[36] ;
 wire \sunrise_digital_top_i.rw_regs[37] ;
 wire \sunrise_digital_top_i.rw_regs[38] ;
 wire \sunrise_digital_top_i.rw_regs[39] ;
 wire \sunrise_digital_top_i.rw_regs[3] ;
 wire \sunrise_digital_top_i.rw_regs[40] ;
 wire \sunrise_digital_top_i.rw_regs[41] ;
 wire \sunrise_digital_top_i.rw_regs[42] ;
 wire \sunrise_digital_top_i.rw_regs[43] ;
 wire \sunrise_digital_top_i.rw_regs[44] ;
 wire \sunrise_digital_top_i.rw_regs[45] ;
 wire \sunrise_digital_top_i.rw_regs[46] ;
 wire \sunrise_digital_top_i.rw_regs[47] ;
 wire \sunrise_digital_top_i.rw_regs[48] ;
 wire \sunrise_digital_top_i.rw_regs[49] ;
 wire \sunrise_digital_top_i.rw_regs[4] ;
 wire \sunrise_digital_top_i.rw_regs[50] ;
 wire \sunrise_digital_top_i.rw_regs[51] ;
 wire \sunrise_digital_top_i.rw_regs[52] ;
 wire \sunrise_digital_top_i.rw_regs[53] ;
 wire \sunrise_digital_top_i.rw_regs[54] ;
 wire \sunrise_digital_top_i.rw_regs[55] ;
 wire \sunrise_digital_top_i.rw_regs[56] ;
 wire \sunrise_digital_top_i.rw_regs[57] ;
 wire \sunrise_digital_top_i.rw_regs[58] ;
 wire \sunrise_digital_top_i.rw_regs[59] ;
 wire \sunrise_digital_top_i.rw_regs[5] ;
 wire \sunrise_digital_top_i.rw_regs[60] ;
 wire \sunrise_digital_top_i.rw_regs[61] ;
 wire \sunrise_digital_top_i.rw_regs[62] ;
 wire \sunrise_digital_top_i.rw_regs[63] ;
 wire \sunrise_digital_top_i.rw_regs[6] ;
 wire \sunrise_digital_top_i.rw_regs[7] ;
 wire \sunrise_digital_top_i.rw_regs[8] ;
 wire \sunrise_digital_top_i.rw_regs[9] ;
 wire \sunrise_digital_top_i.spi_clk_sync ;
 wire \sunrise_digital_top_i.spi_cs_n_sync ;
 wire \sunrise_digital_top_i.spi_mosi_sync ;
 wire \sunrise_digital_top_i.sync_input_prot_sel.data_sync[1] ;
 wire \sunrise_digital_top_i.sync_input_spi_clk.data_sync[1] ;
 wire \sunrise_digital_top_i.sync_input_spi_cpha.data_sync[1] ;
 wire \sunrise_digital_top_i.sync_input_spi_cpol.data_sync[1] ;
 wire \sunrise_digital_top_i.sync_input_spi_cs_n.data_sync[1] ;
 wire \sunrise_digital_top_i.sync_input_spi_mosi.data_sync[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_addr[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_addr[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_addr[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_start ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_stop ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[4] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[5] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[6] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[7] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.pull_sda ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.we ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[10] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[11] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[12] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[17] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[4] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[5] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[6] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[7] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[8] ;
 wire \sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[9] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_sof.data_dly ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_spi_clk.data_dly ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[4] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[5] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[6] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[7] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[4] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[0] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[1] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[2] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[3] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[4] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[5] ;
 wire \sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[6] ;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0592_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[3] ),
    .ZN(_0170_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0593_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[3] ),
    .ZN(_0171_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0594_ (.I(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[17] ),
    .ZN(_0172_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0595_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[2] ),
    .ZN(_0173_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0596_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[3] ),
    .ZN(_0174_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0597_ (.I(\sunrise_digital_top_i.spi_cs_n_sync ),
    .ZN(_0175_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0598_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_sof.data_dly ),
    .ZN(_0176_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0599_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[0] ),
    .ZN(_0177_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0600_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[1] ),
    .ZN(_0178_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0601_ (.I(_0024_),
    .ZN(_0179_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0602_ (.I(_0025_),
    .ZN(_0180_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0603_ (.I(_0026_),
    .ZN(_0181_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0604_ (.I(_0027_),
    .ZN(_0182_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0605_ (.I(_0591_),
    .ZN(_0183_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0606_ (.I(_0016_),
    .ZN(_0184_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0607_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ),
    .ZN(_0185_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0608_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[6] ),
    .ZN(_0186_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0609_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[5] ),
    .ZN(_0187_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0610_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[7] ),
    .ZN(_0188_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0611_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ),
    .ZN(_0189_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0612_ (.I(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[0] ),
    .ZN(_0190_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _0613_ (.I(net47),
    .ZN(_0191_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0614_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ),
    .ZN(_0192_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0615_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[1] ),
    .ZN(_0193_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0616_ (.I(\sunrise_digital_top_i.spi_clk_sync ),
    .ZN(_0194_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0617_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[0] ),
    .ZN(_0195_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0618_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[0] ),
    .ZN(_0196_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0619_ (.I(\sunrise_digital_top_i.rw_regs[33] ),
    .ZN(_0197_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0620_ (.I(\sunrise_digital_top_i.rw_regs[25] ),
    .ZN(_0198_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0621_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[1] ),
    .ZN(_0199_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0622_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[2] ),
    .ZN(_0200_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0623_ (.I(\sunrise_digital_top_i.rw_regs[35] ),
    .ZN(_0201_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0624_ (.I(\sunrise_digital_top_i.rw_regs[27] ),
    .ZN(_0202_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0625_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[3] ),
    .ZN(_0203_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0626_ (.I(\sunrise_digital_top_i.rw_regs[36] ),
    .ZN(_0204_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0627_ (.I(\sunrise_digital_top_i.rw_regs[28] ),
    .ZN(_0205_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0628_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[4] ),
    .ZN(_0206_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0629_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[5] ),
    .ZN(_0207_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0630_ (.I(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[6] ),
    .ZN(_0208_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0631_ (.I(_0030_),
    .ZN(_0209_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _0632_ (.I(net8),
    .ZN(uio_oe[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0633_ (.I(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.pull_sda ),
    .ZN(i2c_sda_oe),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0634_ (.I(spi_miso),
    .ZN(_0210_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0635_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[2] ),
    .A2(_0170_),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ),
    .A4(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[1] ),
    .ZN(_0211_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0636_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[2] ),
    .A2(_0170_),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ),
    .A4(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[1] ),
    .ZN(_0212_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0637_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[3] ),
    .A2(_0212_),
    .B(_0211_),
    .ZN(_0213_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0638_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[0] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[1] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[2] ),
    .ZN(_0214_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0639_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[3] ),
    .A2(_0214_),
    .Z(_0215_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0640_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[3] ),
    .A2(_0214_),
    .ZN(_0216_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0641_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[0] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[1] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[2] ),
    .A4(_0171_),
    .Z(_0217_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0642_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[0] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[1] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[2] ),
    .A4(_0171_),
    .ZN(_0218_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0643_ (.A1(_0213_),
    .A2(net43),
    .A3(_0217_),
    .ZN(_0010_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0644_ (.A1(net69),
    .A2(\sunrise_digital_top_i.spi_cs_n_sync ),
    .ZN(_0219_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0645_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_sof.data_dly ),
    .A2(_0219_),
    .ZN(_0220_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0646_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[1] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[2] ),
    .ZN(_0221_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0647_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[3] ),
    .A2(_0221_),
    .Z(_0222_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0648_ (.I(_0222_),
    .ZN(_0223_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0649_ (.A1(net69),
    .A2(_0222_),
    .Z(_0224_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0650_ (.A1(net70),
    .A2(_0222_),
    .ZN(_0225_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0651_ (.A1(_0220_),
    .A2(_0224_),
    .ZN(_0226_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0652_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[4] ),
    .A2(_0226_),
    .ZN(_0227_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0653_ (.A1(net69),
    .A2(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[2] ),
    .ZN(_0228_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0654_ (.A1(_0172_),
    .A2(_0228_),
    .B(_0227_),
    .ZN(_0015_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0655_ (.A1(\sunrise_digital_top_i.spi_cs_n_sync ),
    .A2(_0176_),
    .ZN(_0229_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0656_ (.A1(net69),
    .A2(_0229_),
    .ZN(_0230_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0657_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[3] ),
    .A2(_0226_),
    .ZN(_0231_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0658_ (.A1(_0177_),
    .A2(_0230_),
    .B(_0231_),
    .ZN(_0014_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0659_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[3] ),
    .A2(_0224_),
    .ZN(_0232_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0660_ (.A1(net69),
    .A2(_0173_),
    .B(_0232_),
    .ZN(_0013_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0661_ (.A1(_0174_),
    .A2(_0221_),
    .Z(_0233_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0662_ (.A1(_0226_),
    .A2(_0233_),
    .ZN(_0234_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0663_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[1] ),
    .A2(_0233_),
    .Z(_0235_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0664_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[1] ),
    .A2(_0233_),
    .ZN(_0236_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0665_ (.A1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[17] ),
    .A2(_0228_),
    .B1(_0234_),
    .B2(_0178_),
    .ZN(_0012_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0666_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[1] ),
    .A2(_0234_),
    .ZN(_0237_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0667_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[4] ),
    .A2(_0224_),
    .ZN(_0238_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0668_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[0] ),
    .A2(_0230_),
    .ZN(_0239_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0669_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[4] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[3] ),
    .B(_0220_),
    .C(_0223_),
    .ZN(_0240_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0670_ (.A1(_0237_),
    .A2(_0238_),
    .A3(_0239_),
    .A4(_0240_),
    .ZN(_0011_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0671_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_stop ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_start ),
    .ZN(_0241_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _0672_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_stop ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_start ),
    .Z(_0242_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0673_ (.A1(_0026_),
    .A2(_0027_),
    .B(_0241_),
    .ZN(_0243_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0674_ (.A1(_0181_),
    .A2(_0182_),
    .B(_0242_),
    .ZN(_0244_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0675_ (.A1(_0179_),
    .A2(_0180_),
    .A3(_0242_),
    .ZN(_0245_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0676_ (.A1(_0024_),
    .A2(_0025_),
    .A3(_0241_),
    .ZN(_0246_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0677_ (.A1(net42),
    .A2(_0245_),
    .ZN(_0247_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0678_ (.A1(_0181_),
    .A2(_0027_),
    .A3(_0242_),
    .ZN(_0248_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0679_ (.A1(_0026_),
    .A2(_0182_),
    .A3(_0241_),
    .ZN(_0249_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0680_ (.A1(_0180_),
    .A2(_0249_),
    .ZN(_0250_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0681_ (.A1(_0025_),
    .A2(_0248_),
    .ZN(_0251_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _0682_ (.A1(_0184_),
    .A2(_0247_),
    .B1(_0251_),
    .B2(_0024_),
    .ZN(_0252_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0683_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[4] ),
    .A4(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ),
    .ZN(_0253_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0684_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[6] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[5] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[7] ),
    .A4(_0253_),
    .ZN(_0254_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0685_ (.A1(_0016_),
    .A2(_0247_),
    .ZN(_0255_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0686_ (.A1(_0016_),
    .A2(_0244_),
    .A3(_0246_),
    .A4(_0254_),
    .ZN(_0256_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0687_ (.A1(_0016_),
    .A2(_0247_),
    .A3(_0254_),
    .Z(_0257_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0688_ (.A1(_0179_),
    .A2(_0025_),
    .A3(_0241_),
    .A4(net42),
    .ZN(_0258_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0689_ (.A1(_0024_),
    .A2(_0248_),
    .ZN(_0259_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0690_ (.A1(_0025_),
    .A2(_0259_),
    .ZN(_0260_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0691_ (.A1(_0024_),
    .A2(_0180_),
    .A3(_0248_),
    .ZN(_0261_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0692_ (.A1(_0258_),
    .A2(_0261_),
    .ZN(_0262_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0693_ (.A1(_0252_),
    .A2(_0256_),
    .A3(_0262_),
    .ZN(_0263_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0694_ (.A1(_0024_),
    .A2(_0025_),
    .B(_0241_),
    .ZN(_0264_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0695_ (.A1(_0179_),
    .A2(_0180_),
    .B(_0242_),
    .ZN(_0265_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0696_ (.A1(_0179_),
    .A2(_0025_),
    .A3(_0242_),
    .ZN(_0266_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0697_ (.A1(_0024_),
    .A2(_0180_),
    .A3(_0241_),
    .ZN(_0267_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0698_ (.A1(_0248_),
    .A2(_0264_),
    .B1(_0266_),
    .B2(_0243_),
    .ZN(_0268_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0699_ (.A1(_0249_),
    .A2(_0265_),
    .B1(_0267_),
    .B2(_0244_),
    .ZN(_0269_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0700_ (.A1(net42),
    .A2(_0264_),
    .ZN(_0270_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _0701_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[3] ),
    .A2(_0591_),
    .A3(_0214_),
    .ZN(_0271_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0702_ (.A1(_0026_),
    .A2(_0182_),
    .A3(_0242_),
    .ZN(_0272_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0703_ (.A1(_0181_),
    .A2(_0027_),
    .A3(_0241_),
    .ZN(_0273_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0704_ (.A1(_0264_),
    .A2(_0272_),
    .ZN(_0274_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0705_ (.A1(_0591_),
    .A2(net43),
    .B(_0274_),
    .ZN(_0275_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0706_ (.A1(_0025_),
    .A2(_0273_),
    .ZN(_0276_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0707_ (.A1(_0180_),
    .A2(_0272_),
    .ZN(_0277_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0708_ (.A1(_0266_),
    .A2(_0272_),
    .ZN(_0278_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0709_ (.I0(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ),
    .I1(net43),
    .S(_0218_),
    .Z(_0279_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0710_ (.A1(_0242_),
    .A2(_0270_),
    .B1(_0278_),
    .B2(_0279_),
    .ZN(_0280_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0711_ (.A1(_0275_),
    .A2(_0280_),
    .ZN(_0281_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _0712_ (.A1(net43),
    .A2(_0263_),
    .B1(_0268_),
    .B2(_0217_),
    .C(_0281_),
    .ZN(_0282_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0713_ (.A1(_0164_),
    .A2(_0162_),
    .A3(_0169_),
    .A4(_0167_),
    .Z(_0283_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0714_ (.A1(net15),
    .A2(_0283_),
    .ZN(_0284_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0715_ (.A1(_0591_),
    .A2(_0261_),
    .ZN(_0285_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0716_ (.A1(_0252_),
    .A2(_0285_),
    .B(net43),
    .ZN(_0286_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0717_ (.A1(_0257_),
    .A2(_0278_),
    .ZN(_0287_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0718_ (.A1(_0189_),
    .A2(_0278_),
    .ZN(_0288_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0719_ (.A1(_0215_),
    .A2(_0287_),
    .A3(_0288_),
    .ZN(_0289_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0720_ (.A1(_0218_),
    .A2(_0249_),
    .A3(_0265_),
    .ZN(_0290_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0721_ (.A1(_0591_),
    .A2(net43),
    .A3(_0260_),
    .ZN(_0291_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0722_ (.I(_0291_),
    .ZN(_0023_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0723_ (.A1(_0290_),
    .A2(_0023_),
    .ZN(_0292_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0724_ (.A1(_0284_),
    .A2(_0286_),
    .A3(_0289_),
    .A4(_0292_),
    .ZN(_0019_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0725_ (.A1(_0162_),
    .A2(net15),
    .ZN(_0293_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0726_ (.A1(_0286_),
    .A2(_0293_),
    .ZN(_0001_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0727_ (.A1(_0258_),
    .A2(_0271_),
    .Z(_0294_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0728_ (.A1(_0289_),
    .A2(_0294_),
    .Z(_0295_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0729_ (.A1(_0217_),
    .A2(_0243_),
    .A3(_0266_),
    .ZN(_0296_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0730_ (.A1(_0168_),
    .A2(net15),
    .ZN(_0297_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0731_ (.A1(_0164_),
    .A2(_0169_),
    .A3(_0163_),
    .A4(_0168_),
    .Z(_0298_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0732_ (.A1(net15),
    .A2(_0298_),
    .ZN(_0299_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0733_ (.A1(_0291_),
    .A2(_0295_),
    .A3(_0296_),
    .A4(_0299_),
    .ZN(_0018_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0734_ (.A1(_0024_),
    .A2(_0250_),
    .ZN(_0300_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0735_ (.A1(_0161_),
    .A2(net15),
    .ZN(_0301_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0736_ (.A1(_0300_),
    .A2(_0301_),
    .ZN(_0000_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0737_ (.A1(_0169_),
    .A2(_0167_),
    .A3(_0168_),
    .A4(_0165_),
    .Z(_0302_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0738_ (.A1(_0166_),
    .A2(_0302_),
    .B(net15),
    .ZN(_0303_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0739_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ),
    .A2(_0257_),
    .ZN(_0304_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0740_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ),
    .A2(_0257_),
    .B1(_0258_),
    .B2(_0591_),
    .ZN(_0305_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0741_ (.A1(net43),
    .A2(_0305_),
    .B(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_start ),
    .ZN(_0306_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0742_ (.A1(_0271_),
    .A2(_0274_),
    .ZN(_0307_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0743_ (.A1(_0290_),
    .A2(_0307_),
    .ZN(_0308_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0744_ (.A1(_0295_),
    .A2(_0303_),
    .A3(_0306_),
    .A4(_0308_),
    .ZN(_0017_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0745_ (.A1(_0169_),
    .A2(net15),
    .ZN(_0309_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0746_ (.A1(_0289_),
    .A2(_0309_),
    .ZN(_0008_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0747_ (.A1(_0294_),
    .A2(_0297_),
    .ZN(_0007_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0748_ (.A1(_0167_),
    .A2(net15),
    .B(_0290_),
    .ZN(_0310_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0749_ (.I(_0310_),
    .ZN(_0006_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0750_ (.A1(_0166_),
    .A2(net15),
    .B(_0307_),
    .ZN(_0311_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0751_ (.I(_0311_),
    .ZN(_0005_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0752_ (.A1(_0212_),
    .A2(_0216_),
    .ZN(_0312_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0753_ (.A1(_0195_),
    .A2(_0211_),
    .A3(_0312_),
    .B(_0218_),
    .ZN(_0009_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0754_ (.A1(_0163_),
    .A2(net15),
    .ZN(_0313_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0755_ (.A1(_0296_),
    .A2(_0313_),
    .ZN(_0002_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0756_ (.A1(_0164_),
    .A2(_0282_),
    .ZN(_0314_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0757_ (.A1(_0291_),
    .A2(_0314_),
    .ZN(_0003_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0758_ (.A1(_0300_),
    .A2(_0301_),
    .A3(_0311_),
    .ZN(_0020_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0759_ (.A1(_0165_),
    .A2(_0282_),
    .ZN(_0315_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0760_ (.A1(_0306_),
    .A2(_0315_),
    .ZN(_0004_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0761_ (.A1(_0195_),
    .A2(_0212_),
    .ZN(_0022_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0762_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[3] ),
    .A2(net43),
    .Z(_0021_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0763_ (.A1(net69),
    .A2(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_spi_clk.data_dly ),
    .ZN(_0316_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0764_ (.A1(net69),
    .A2(_0194_),
    .B(_0316_),
    .ZN(_0031_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0765_ (.A1(net69),
    .A2(_0176_),
    .B(_0219_),
    .ZN(_0032_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0766_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[0] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[1] ),
    .S(_0238_),
    .Z(_0033_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0767_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[1] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[2] ),
    .S(_0238_),
    .Z(_0034_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0768_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[2] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[3] ),
    .S(_0238_),
    .Z(_0035_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0769_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[3] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[4] ),
    .S(_0238_),
    .Z(_0036_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0770_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[4] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[5] ),
    .S(_0238_),
    .Z(_0037_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0771_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[5] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[6] ),
    .S(_0238_),
    .Z(_0038_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0772_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[6] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[7] ),
    .S(_0238_),
    .Z(_0039_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0773_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[7] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[8] ),
    .S(_0238_),
    .Z(_0040_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0774_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[0] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[9] ),
    .S(_0232_),
    .Z(_0041_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0775_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[1] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[10] ),
    .S(_0232_),
    .Z(_0042_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0776_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[2] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[11] ),
    .S(_0232_),
    .Z(_0043_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0777_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[3] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[12] ),
    .S(_0232_),
    .Z(_0044_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0778_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[7] ),
    .A2(_0232_),
    .ZN(_0317_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0779_ (.A1(_0172_),
    .A2(_0232_),
    .B(_0317_),
    .ZN(_0045_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0780_ (.A1(net70),
    .A2(_0190_),
    .B1(_0238_),
    .B2(_0172_),
    .ZN(_0046_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _0781_ (.A1(\sunrise_digital_top_i.cpha_sync ),
    .A2(\sunrise_digital_top_i.cpol_sync ),
    .Z(_0318_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0782_ (.A1(_0175_),
    .A2(_0194_),
    .A3(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_spi_clk.data_dly ),
    .ZN(_0319_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0783_ (.A1(_0318_),
    .A2(_0319_),
    .ZN(_0320_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0784_ (.A1(\sunrise_digital_top_i.spi_cs_n_sync ),
    .A2(_0194_),
    .A3(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_spi_clk.data_dly ),
    .ZN(_0321_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _0785_ (.A1(_0318_),
    .A2(_0321_),
    .B(_0320_),
    .C(net69),
    .ZN(_0322_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0786_ (.A1(_0225_),
    .A2(net37),
    .ZN(_0323_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0787_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ),
    .A2(_0323_),
    .ZN(_0324_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0788_ (.A1(_0222_),
    .A2(net37),
    .ZN(_0325_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0789_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ),
    .A2(_0325_),
    .B(_0324_),
    .ZN(_0326_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0790_ (.I(_0326_),
    .ZN(_0047_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0791_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[1] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ),
    .A3(_0323_),
    .ZN(_0327_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0792_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[1] ),
    .A2(_0324_),
    .ZN(_0048_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0793_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[1] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[2] ),
    .ZN(_0328_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0794_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[2] ),
    .A2(_0327_),
    .ZN(_0049_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0795_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[3] ),
    .A2(_0328_),
    .Z(_0329_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0796_ (.A1(_0222_),
    .A2(net37),
    .A3(_0329_),
    .B1(_0323_),
    .B2(_0174_),
    .ZN(_0050_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0797_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.we ),
    .A2(_0191_),
    .B(net68),
    .ZN(_0330_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0798_ (.A1(_0190_),
    .A2(_0191_),
    .B(_0330_),
    .ZN(_0331_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0799_ (.A1(net46),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[10] ),
    .ZN(_0332_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0800_ (.I0(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[10] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[1] ),
    .S(net48),
    .Z(_0333_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0801_ (.A1(net46),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[9] ),
    .ZN(_0334_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0802_ (.I0(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[9] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ),
    .S(net46),
    .Z(_0335_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0803_ (.A1(_0333_),
    .A2(net45),
    .Z(_0336_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0804_ (.A1(_0333_),
    .A2(net45),
    .ZN(_0337_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0805_ (.A1(net47),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[2] ),
    .Z(_0338_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0806_ (.A1(_0191_),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[11] ),
    .B(_0338_),
    .ZN(_0339_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0807_ (.I0(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[11] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[2] ),
    .S(net47),
    .Z(_0340_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0808_ (.A1(_0333_),
    .A2(net45),
    .A3(net44),
    .Z(_0341_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0809_ (.A1(_0331_),
    .A2(_0341_),
    .ZN(_0342_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0810_ (.A1(_0189_),
    .A2(net46),
    .ZN(_0343_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0811_ (.A1(net46),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[1] ),
    .B(_0343_),
    .ZN(_0344_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0812_ (.A1(\sunrise_digital_top_i.rw_regs[56] ),
    .A2(net35),
    .ZN(_0345_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0813_ (.A1(net35),
    .A2(_0344_),
    .B(_0345_),
    .ZN(_0051_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0814_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .A2(net47),
    .Z(_0346_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0815_ (.A1(_0191_),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[2] ),
    .B(_0346_),
    .ZN(_0347_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0816_ (.I0(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[2] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .S(net48),
    .Z(_0348_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0817_ (.A1(\sunrise_digital_top_i.rw_regs[57] ),
    .A2(net35),
    .ZN(_0349_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0818_ (.A1(net36),
    .A2(_0347_),
    .B(_0349_),
    .ZN(_0052_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0819_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ),
    .A2(net47),
    .Z(_0350_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0820_ (.A1(_0191_),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[3] ),
    .B(_0350_),
    .ZN(_0351_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0821_ (.A1(\sunrise_digital_top_i.rw_regs[58] ),
    .A2(net35),
    .ZN(_0352_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0822_ (.A1(net35),
    .A2(_0351_),
    .B(_0352_),
    .ZN(_0053_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0823_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ),
    .A2(net47),
    .ZN(_0353_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0824_ (.A1(_0191_),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[4] ),
    .ZN(_0354_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0825_ (.A1(_0353_),
    .A2(_0354_),
    .Z(_0355_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0826_ (.A1(_0353_),
    .A2(_0354_),
    .ZN(_0356_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0827_ (.A1(\sunrise_digital_top_i.rw_regs[59] ),
    .A2(net36),
    .ZN(_0357_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0828_ (.A1(net36),
    .A2(_0355_),
    .B(_0357_),
    .ZN(_0054_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0829_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[4] ),
    .A2(net47),
    .Z(_0358_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0830_ (.A1(_0191_),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[5] ),
    .B(_0358_),
    .ZN(_0359_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0831_ (.A1(\sunrise_digital_top_i.rw_regs[60] ),
    .A2(net36),
    .ZN(_0360_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0832_ (.A1(net36),
    .A2(_0359_),
    .B(_0360_),
    .ZN(_0055_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0833_ (.A1(_0187_),
    .A2(net46),
    .ZN(_0361_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0834_ (.A1(net47),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[6] ),
    .B(_0361_),
    .ZN(_0362_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0835_ (.A1(\sunrise_digital_top_i.rw_regs[61] ),
    .A2(net36),
    .ZN(_0363_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0836_ (.A1(net35),
    .A2(_0362_),
    .B(_0363_),
    .ZN(_0056_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0837_ (.A1(_0186_),
    .A2(net46),
    .ZN(_0364_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0838_ (.A1(net46),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[7] ),
    .B(_0364_),
    .ZN(_0365_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0839_ (.A1(\sunrise_digital_top_i.rw_regs[62] ),
    .A2(net35),
    .ZN(_0366_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0840_ (.A1(net35),
    .A2(_0365_),
    .B(_0366_),
    .ZN(_0057_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0841_ (.A1(_0188_),
    .A2(net46),
    .ZN(_0367_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0842_ (.A1(net46),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[8] ),
    .B(_0367_),
    .ZN(_0368_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0843_ (.A1(\sunrise_digital_top_i.rw_regs[63] ),
    .A2(net35),
    .ZN(_0369_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0844_ (.A1(net35),
    .A2(_0368_),
    .B(_0369_),
    .ZN(_0058_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0845_ (.A1(net68),
    .A2(_0235_),
    .ZN(_0370_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0846_ (.A1(_0318_),
    .A2(_0321_),
    .ZN(_0371_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0847_ (.A1(_0318_),
    .A2(_0319_),
    .B(_0371_),
    .ZN(_0372_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0848_ (.A1(_0235_),
    .A2(_0372_),
    .B(net69),
    .ZN(_0373_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0849_ (.A1(_0230_),
    .A2(_0373_),
    .ZN(_0374_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0850_ (.A1(_0337_),
    .A2(net44),
    .ZN(_0375_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0851_ (.A1(net47),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[3] ),
    .Z(_0376_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _0852_ (.A1(_0191_),
    .A2(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[12] ),
    .B(_0376_),
    .ZN(_0377_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0853_ (.I0(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[12] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[3] ),
    .S(net47),
    .Z(_0378_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0854_ (.A1(_0375_),
    .A2(net41),
    .ZN(_0379_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0855_ (.A1(net45),
    .A2(_0339_),
    .B(_0379_),
    .ZN(_0380_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0856_ (.A1(_0333_),
    .A2(net45),
    .ZN(_0381_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0857_ (.A1(_0333_),
    .A2(net45),
    .Z(_0382_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0858_ (.A1(net44),
    .A2(_0382_),
    .ZN(_0383_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0859_ (.A1(_0339_),
    .A2(_0381_),
    .ZN(_0384_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _0860_ (.A1(net98),
    .A2(_0193_),
    .B(net45),
    .C(_0332_),
    .ZN(_0385_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0861_ (.A1(net44),
    .A2(net94),
    .Z(_0386_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0862_ (.A1(_0339_),
    .A2(_0385_),
    .Z(_0387_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _0863_ (.A1(net97),
    .A2(_0192_),
    .B(_0333_),
    .C(_0334_),
    .ZN(_0388_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _0864_ (.A1(_0339_),
    .A2(_0388_),
    .Z(_0389_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _0865_ (.A1(net44),
    .A2(_0388_),
    .Z(_0390_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0866_ (.A1(\sunrise_digital_top_i.rw_regs[56] ),
    .A2(_0341_),
    .B1(_0381_),
    .B2(\sunrise_digital_top_i.rw_regs[32] ),
    .C1(_0390_),
    .C2(\sunrise_digital_top_i.rw_regs[40] ),
    .ZN(_0391_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0867_ (.A1(\sunrise_digital_top_i.rw_regs[48] ),
    .A2(_0386_),
    .B1(_0389_),
    .B2(\sunrise_digital_top_i.rw_regs[8] ),
    .ZN(_0392_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0868_ (.A1(\sunrise_digital_top_i.rw_regs[24] ),
    .A2(_0375_),
    .B1(_0387_),
    .B2(\sunrise_digital_top_i.rw_regs[16] ),
    .ZN(_0393_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0869_ (.A1(_0391_),
    .A2(_0392_),
    .A3(_0393_),
    .Z(_0394_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0870_ (.A1(\sunrise_digital_top_i.rw_regs[0] ),
    .A2(net39),
    .ZN(_0395_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0871_ (.A1(net39),
    .A2(_0394_),
    .B(_0395_),
    .C(net41),
    .ZN(_0396_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0872_ (.A1(_0380_),
    .A2(_0396_),
    .ZN(_0397_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0873_ (.A1(_0229_),
    .A2(_0370_),
    .A3(_0397_),
    .B1(_0374_),
    .B2(_0196_),
    .ZN(_0059_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0874_ (.A1(_0336_),
    .A2(_0381_),
    .B(net44),
    .ZN(_0398_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0875_ (.A1(net45),
    .A2(_0340_),
    .B(_0378_),
    .C(_0398_),
    .ZN(_0399_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0876_ (.A1(\sunrise_digital_top_i.rw_regs[57] ),
    .A2(_0341_),
    .B1(_0386_),
    .B2(\sunrise_digital_top_i.rw_regs[49] ),
    .C1(_0390_),
    .C2(\sunrise_digital_top_i.rw_regs[41] ),
    .ZN(_0400_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0877_ (.A1(_0198_),
    .A2(_0337_),
    .A3(net44),
    .B1(_0382_),
    .B2(_0197_),
    .ZN(_0401_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0878_ (.A1(\sunrise_digital_top_i.rw_regs[17] ),
    .A2(net93),
    .B1(_0389_),
    .B2(\sunrise_digital_top_i.rw_regs[9] ),
    .C(_0401_),
    .ZN(_0402_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0879_ (.A1(net34),
    .A2(_0402_),
    .B(net40),
    .ZN(_0403_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0880_ (.A1(\sunrise_digital_top_i.rw_regs[1] ),
    .A2(net39),
    .ZN(_0404_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0881_ (.A1(net41),
    .A2(_0404_),
    .ZN(_0405_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0882_ (.A1(_0403_),
    .A2(_0405_),
    .B(_0399_),
    .ZN(_0406_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0883_ (.A1(_0229_),
    .A2(_0373_),
    .Z(_0407_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0884_ (.I0(_0196_),
    .I1(_0406_),
    .S(_0235_),
    .Z(_0408_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0885_ (.A1(_0199_),
    .A2(_0374_),
    .B1(_0407_),
    .B2(_0408_),
    .ZN(_0060_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0886_ (.A1(\sunrise_digital_top_i.rw_regs[26] ),
    .A2(_0375_),
    .B1(net93),
    .B2(\sunrise_digital_top_i.rw_regs[18] ),
    .C1(_0390_),
    .C2(\sunrise_digital_top_i.rw_regs[42] ),
    .ZN(_0409_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0887_ (.A1(\sunrise_digital_top_i.rw_regs[10] ),
    .A2(_0339_),
    .A3(_0388_),
    .ZN(_0410_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0888_ (.A1(\sunrise_digital_top_i.rw_regs[34] ),
    .A2(_0381_),
    .ZN(_0411_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0889_ (.A1(\sunrise_digital_top_i.rw_regs[50] ),
    .A2(net44),
    .A3(net94),
    .ZN(_0412_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0890_ (.A1(\sunrise_digital_top_i.rw_regs[58] ),
    .A2(_0341_),
    .ZN(_0413_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0891_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0412_),
    .A4(_0413_),
    .Z(_0414_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0892_ (.A1(_0409_),
    .A2(_0414_),
    .B(net39),
    .ZN(_0415_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0893_ (.A1(\sunrise_digital_top_i.rw_regs[2] ),
    .A2(net39),
    .ZN(_0416_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0894_ (.A1(net41),
    .A2(_0416_),
    .ZN(_0417_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0895_ (.A1(_0415_),
    .A2(_0417_),
    .B(_0380_),
    .ZN(_0418_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0896_ (.I0(_0199_),
    .I1(_0418_),
    .S(_0235_),
    .Z(_0419_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0897_ (.A1(_0200_),
    .A2(_0374_),
    .B1(_0407_),
    .B2(_0419_),
    .ZN(_0061_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0898_ (.A1(\sunrise_digital_top_i.rw_regs[59] ),
    .A2(_0341_),
    .B1(_0387_),
    .B2(\sunrise_digital_top_i.rw_regs[19] ),
    .C1(_0390_),
    .C2(\sunrise_digital_top_i.rw_regs[43] ),
    .ZN(_0420_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0899_ (.A1(_0202_),
    .A2(_0337_),
    .A3(_0340_),
    .B1(_0382_),
    .B2(_0201_),
    .ZN(_0421_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0900_ (.A1(\sunrise_digital_top_i.rw_regs[51] ),
    .A2(_0386_),
    .B1(_0389_),
    .B2(\sunrise_digital_top_i.rw_regs[11] ),
    .C(net38),
    .ZN(_0422_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0901_ (.A1(net33),
    .A2(_0422_),
    .B(net40),
    .ZN(_0423_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0902_ (.A1(\sunrise_digital_top_i.rw_regs[3] ),
    .A2(net39),
    .ZN(_0424_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0903_ (.A1(net41),
    .A2(_0424_),
    .ZN(_0425_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0904_ (.A1(_0423_),
    .A2(_0425_),
    .B(_0399_),
    .ZN(_0426_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0905_ (.I0(_0200_),
    .I1(_0426_),
    .S(_0235_),
    .Z(_0427_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0906_ (.A1(_0203_),
    .A2(_0374_),
    .B1(_0407_),
    .B2(_0427_),
    .ZN(_0062_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0907_ (.A1(\sunrise_digital_top_i.rw_regs[52] ),
    .A2(_0386_),
    .B1(_0389_),
    .B2(\sunrise_digital_top_i.rw_regs[12] ),
    .C1(_0390_),
    .C2(\sunrise_digital_top_i.rw_regs[44] ),
    .ZN(_0428_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0908_ (.A1(_0205_),
    .A2(_0337_),
    .A3(net44),
    .B1(_0382_),
    .B2(_0204_),
    .ZN(_0429_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0909_ (.A1(\sunrise_digital_top_i.rw_regs[60] ),
    .A2(_0341_),
    .B1(net93),
    .B2(\sunrise_digital_top_i.rw_regs[20] ),
    .C(_0429_),
    .ZN(_0430_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0910_ (.A1(net32),
    .A2(_0430_),
    .B(net40),
    .ZN(_0431_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0911_ (.A1(\sunrise_digital_top_i.rw_regs[4] ),
    .A2(net40),
    .ZN(_0432_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0912_ (.A1(_0377_),
    .A2(_0432_),
    .ZN(_0433_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0913_ (.A1(net45),
    .A2(_0339_),
    .B(net41),
    .ZN(_0434_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0914_ (.A1(_0398_),
    .A2(_0434_),
    .ZN(_0435_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0915_ (.A1(_0431_),
    .A2(_0433_),
    .B(_0435_),
    .ZN(_0436_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0916_ (.I0(_0203_),
    .I1(_0436_),
    .S(_0235_),
    .Z(_0437_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _0917_ (.A1(_0206_),
    .A2(_0374_),
    .B1(_0407_),
    .B2(_0437_),
    .ZN(_0063_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0918_ (.A1(\sunrise_digital_top_i.rw_regs[53] ),
    .A2(_0386_),
    .B1(_0390_),
    .B2(\sunrise_digital_top_i.rw_regs[45] ),
    .C1(\sunrise_digital_top_i.rw_regs[29] ),
    .C2(_0375_),
    .ZN(_0438_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0919_ (.A1(\sunrise_digital_top_i.rw_regs[61] ),
    .A2(_0341_),
    .B1(_0381_),
    .B2(\sunrise_digital_top_i.rw_regs[37] ),
    .C(net39),
    .ZN(_0439_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0920_ (.A1(\sunrise_digital_top_i.rw_regs[21] ),
    .A2(_0387_),
    .B1(_0389_),
    .B2(\sunrise_digital_top_i.rw_regs[13] ),
    .ZN(_0440_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0921_ (.A1(_0438_),
    .A2(_0439_),
    .A3(_0440_),
    .Z(_0441_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0922_ (.A1(\sunrise_digital_top_i.rw_regs[5] ),
    .A2(_0384_),
    .B(_0377_),
    .ZN(_0442_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0923_ (.A1(_0335_),
    .A2(_0377_),
    .A3(net39),
    .B1(_0441_),
    .B2(_0442_),
    .ZN(_0443_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0924_ (.A1(_0236_),
    .A2(net14),
    .ZN(_0444_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0925_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[4] ),
    .A2(_0235_),
    .ZN(_0445_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0926_ (.A1(_0407_),
    .A2(_0444_),
    .A3(_0445_),
    .B1(_0374_),
    .B2(_0207_),
    .ZN(_0064_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0927_ (.A1(\sunrise_digital_top_i.rw_regs[62] ),
    .A2(_0341_),
    .B1(_0381_),
    .B2(\sunrise_digital_top_i.rw_regs[38] ),
    .C(net39),
    .ZN(_0446_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0928_ (.A1(\sunrise_digital_top_i.rw_regs[30] ),
    .A2(_0375_),
    .B1(_0387_),
    .B2(\sunrise_digital_top_i.rw_regs[22] ),
    .C1(_0390_),
    .C2(\sunrise_digital_top_i.rw_regs[46] ),
    .ZN(_0447_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0929_ (.A1(\sunrise_digital_top_i.rw_regs[54] ),
    .A2(_0386_),
    .B1(_0389_),
    .B2(\sunrise_digital_top_i.rw_regs[14] ),
    .ZN(_0448_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _0930_ (.A1(_0446_),
    .A2(_0447_),
    .A3(_0448_),
    .Z(_0449_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0931_ (.A1(\sunrise_digital_top_i.rw_regs[6] ),
    .A2(_0384_),
    .B(net41),
    .ZN(_0450_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _0932_ (.A1(net41),
    .A2(net96),
    .A3(_0388_),
    .B1(_0449_),
    .B2(_0450_),
    .ZN(_0451_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0933_ (.A1(_0236_),
    .A2(net13),
    .ZN(_0452_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0934_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[5] ),
    .A2(_0235_),
    .ZN(_0453_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0935_ (.A1(_0407_),
    .A2(_0452_),
    .A3(_0453_),
    .B1(_0374_),
    .B2(_0208_),
    .ZN(_0065_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0936_ (.A1(\sunrise_digital_top_i.rw_regs[31] ),
    .A2(_0375_),
    .B1(_0387_),
    .B2(\sunrise_digital_top_i.rw_regs[23] ),
    .C1(_0389_),
    .C2(\sunrise_digital_top_i.rw_regs[15] ),
    .ZN(_0454_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0937_ (.A1(\sunrise_digital_top_i.rw_regs[63] ),
    .A2(_0341_),
    .B1(_0390_),
    .B2(\sunrise_digital_top_i.rw_regs[47] ),
    .ZN(_0455_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0938_ (.A1(\sunrise_digital_top_i.rw_regs[39] ),
    .A2(_0381_),
    .B1(_0386_),
    .B2(\sunrise_digital_top_i.rw_regs[55] ),
    .C(net39),
    .ZN(_0456_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0939_ (.A1(_0454_),
    .A2(_0455_),
    .A3(_0456_),
    .Z(_0457_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0940_ (.A1(\sunrise_digital_top_i.rw_regs[7] ),
    .A2(_0384_),
    .B(net41),
    .ZN(_0458_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _0941_ (.A1(net45),
    .A2(net41),
    .B1(_0457_),
    .B2(_0458_),
    .ZN(_0459_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0942_ (.A1(_0236_),
    .A2(_0459_),
    .ZN(_0460_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0943_ (.A1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[6] ),
    .A2(_0235_),
    .ZN(_0461_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0944_ (.A1(_0407_),
    .A2(_0460_),
    .A3(_0461_),
    .B1(_0374_),
    .B2(_0210_),
    .ZN(_0066_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0945_ (.I0(\sunrise_digital_top_i.spi_mosi_sync ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[0] ),
    .S(net37),
    .Z(_0067_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0946_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[0] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[1] ),
    .S(net37),
    .Z(_0068_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0947_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[1] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[2] ),
    .S(net37),
    .Z(_0069_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0948_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[2] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[3] ),
    .S(net37),
    .Z(_0070_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0949_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[3] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[4] ),
    .S(net37),
    .Z(_0071_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0950_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[4] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[5] ),
    .S(net37),
    .Z(_0072_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0951_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[5] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[6] ),
    .S(net37),
    .Z(_0073_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0952_ (.I0(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[6] ),
    .I1(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[7] ),
    .S(_0322_),
    .Z(_0074_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0953_ (.A1(_0256_),
    .A2(_0276_),
    .B(_0216_),
    .ZN(_0462_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0954_ (.A1(_0184_),
    .A2(net42),
    .A3(_0245_),
    .A4(_0254_),
    .ZN(_0463_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _0955_ (.A1(_0184_),
    .A2(_0244_),
    .A3(_0246_),
    .B1(_0265_),
    .B2(_0271_),
    .B3(_0273_),
    .ZN(_0464_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0956_ (.A1(_0218_),
    .A2(_0269_),
    .B(_0464_),
    .ZN(_0465_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0957_ (.A1(_0247_),
    .A2(_0268_),
    .A3(_0277_),
    .ZN(_0466_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0958_ (.A1(_0247_),
    .A2(_0268_),
    .A3(_0270_),
    .A4(_0277_),
    .ZN(_0467_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0959_ (.A1(_0462_),
    .A2(_0463_),
    .A3(_0465_),
    .A4(_0467_),
    .ZN(_0468_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0960_ (.A1(_0304_),
    .A2(_0468_),
    .Z(_0469_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0961_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .A2(net12),
    .ZN(_0470_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0962_ (.A1(_0268_),
    .A2(_0274_),
    .ZN(_0471_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0963_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ),
    .A2(net30),
    .ZN(_0472_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0964_ (.A1(_0406_),
    .A2(_0472_),
    .Z(_0473_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0965_ (.A1(_0288_),
    .A2(_0466_),
    .ZN(_0474_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0966_ (.A1(net12),
    .A2(_0473_),
    .A3(_0474_),
    .B(_0470_),
    .ZN(_0075_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0967_ (.A1(_0189_),
    .A2(_0247_),
    .B(_0278_),
    .ZN(_0475_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0968_ (.I(_0475_),
    .ZN(_0476_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0969_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .A2(net30),
    .ZN(_0477_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0970_ (.A1(_0418_),
    .A2(_0476_),
    .B(_0477_),
    .ZN(_0478_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0971_ (.I0(_0478_),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ),
    .S(net12),
    .Z(_0076_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0972_ (.A1(_0426_),
    .A2(_0476_),
    .Z(_0479_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0973_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ),
    .A2(net30),
    .B(net12),
    .ZN(_0480_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0974_ (.A1(_0185_),
    .A2(net12),
    .B1(_0479_),
    .B2(_0480_),
    .ZN(_0077_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0975_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ),
    .A2(net30),
    .ZN(_0481_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0976_ (.A1(_0436_),
    .A2(_0476_),
    .B(_0481_),
    .ZN(_0482_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0977_ (.I0(_0482_),
    .I1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[4] ),
    .S(net12),
    .Z(_0078_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0978_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[4] ),
    .A2(_0471_),
    .B1(_0475_),
    .B2(_0443_),
    .C(_0469_),
    .ZN(_0483_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0979_ (.A1(_0187_),
    .A2(_0469_),
    .B(_0483_),
    .ZN(_0079_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0980_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[5] ),
    .A2(_0471_),
    .B1(_0475_),
    .B2(_0451_),
    .C(net12),
    .ZN(_0484_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0981_ (.A1(_0186_),
    .A2(net12),
    .B(_0484_),
    .ZN(_0080_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0982_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[6] ),
    .A2(_0471_),
    .B1(_0475_),
    .B2(_0459_),
    .C(net12),
    .ZN(_0485_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0983_ (.A1(_0188_),
    .A2(net12),
    .B(_0485_),
    .ZN(_0081_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0984_ (.A1(_0180_),
    .A2(_0182_),
    .B(_0242_),
    .ZN(_0486_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0985_ (.A1(_0258_),
    .A2(_0274_),
    .A3(_0486_),
    .ZN(_0487_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0986_ (.A1(_0024_),
    .A2(_0251_),
    .B(_0247_),
    .ZN(_0488_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0987_ (.A1(_0487_),
    .A2(_0488_),
    .B(_0463_),
    .ZN(_0489_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0988_ (.A1(net43),
    .A2(_0488_),
    .ZN(_0490_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0989_ (.A1(net43),
    .A2(_0488_),
    .B(_0487_),
    .ZN(_0491_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0990_ (.A1(_0188_),
    .A2(_0275_),
    .B(_0491_),
    .ZN(_0492_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0991_ (.A1(i2c_sda_oe),
    .A2(_0489_),
    .B1(_0492_),
    .B2(_0463_),
    .ZN(_0082_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0992_ (.A1(_0216_),
    .A2(_0247_),
    .A3(_0254_),
    .ZN(_0493_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0993_ (.A1(_0016_),
    .A2(_0493_),
    .B(_0270_),
    .ZN(_0494_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0994_ (.I(_0494_),
    .ZN(_0083_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _0995_ (.A1(_0300_),
    .A2(_0490_),
    .B(_0255_),
    .ZN(_0495_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0996_ (.A1(_0192_),
    .A2(_0250_),
    .B1(_0300_),
    .B2(_0490_),
    .C(_0255_),
    .ZN(_0496_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0997_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ),
    .A2(_0251_),
    .B(_0495_),
    .ZN(_0497_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0998_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ),
    .A2(_0251_),
    .ZN(_0498_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0999_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ),
    .A2(_0495_),
    .ZN(_0499_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1000_ (.A1(_0496_),
    .A2(_0498_),
    .B(_0499_),
    .ZN(_0084_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1001_ (.A1(_0192_),
    .A2(_0193_),
    .B(_0250_),
    .ZN(_0500_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1002_ (.A1(_0495_),
    .A2(_0500_),
    .Z(_0501_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1003_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .A2(_0251_),
    .ZN(_0502_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1004_ (.A1(_0193_),
    .A2(_0497_),
    .B1(_0501_),
    .B2(_0502_),
    .ZN(_0085_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1005_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ),
    .A2(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[1] ),
    .A3(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[2] ),
    .ZN(_0503_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1006_ (.A1(_0251_),
    .A2(_0503_),
    .Z(_0504_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1007_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ),
    .A2(_0250_),
    .B(_0504_),
    .ZN(_0505_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1008_ (.A1(_0495_),
    .A2(_0500_),
    .B(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[2] ),
    .ZN(_0506_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1009_ (.A1(_0495_),
    .A2(_0505_),
    .B(_0506_),
    .ZN(_0086_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1010_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[3] ),
    .A2(_0503_),
    .Z(_0507_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1011_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ),
    .A2(_0251_),
    .ZN(_0508_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1012_ (.A1(_0251_),
    .A2(_0507_),
    .B(_0508_),
    .ZN(_0509_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1013_ (.I0(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[3] ),
    .I1(_0509_),
    .S(_0495_),
    .Z(_0087_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1014_ (.I0(\sunrise_digital_top_i.spi_mosi_sync ),
    .I1(\sunrise_digital_top_i.sync_input_spi_mosi.data_sync[1] ),
    .S(net68),
    .Z(_0088_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1015_ (.A1(_0380_),
    .A2(_0396_),
    .A3(_0475_),
    .ZN(_0510_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1016_ (.A1(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ),
    .A2(_0269_),
    .B(_0468_),
    .ZN(_0511_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1017_ (.A1(_0189_),
    .A2(_0468_),
    .B1(_0510_),
    .B2(_0511_),
    .ZN(_0089_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1018_ (.A1(_0331_),
    .A2(net44),
    .A3(_0381_),
    .ZN(_0512_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1019_ (.A1(\sunrise_digital_top_i.rw_regs[32] ),
    .A2(net28),
    .ZN(_0513_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1020_ (.A1(_0344_),
    .A2(net28),
    .B(_0513_),
    .ZN(_0090_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1021_ (.A1(\sunrise_digital_top_i.rw_regs[33] ),
    .A2(net29),
    .ZN(_0514_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1022_ (.A1(_0347_),
    .A2(net29),
    .B(_0514_),
    .ZN(_0091_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1023_ (.A1(\sunrise_digital_top_i.rw_regs[34] ),
    .A2(net28),
    .ZN(_0515_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1024_ (.A1(_0351_),
    .A2(net28),
    .B(_0515_),
    .ZN(_0092_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1025_ (.A1(\sunrise_digital_top_i.rw_regs[35] ),
    .A2(net29),
    .ZN(_0516_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1026_ (.A1(_0355_),
    .A2(net29),
    .B(_0516_),
    .ZN(_0093_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1027_ (.A1(\sunrise_digital_top_i.rw_regs[36] ),
    .A2(net29),
    .ZN(_0517_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1028_ (.A1(_0359_),
    .A2(net29),
    .B(_0517_),
    .ZN(_0094_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1029_ (.A1(\sunrise_digital_top_i.rw_regs[37] ),
    .A2(net28),
    .ZN(_0518_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1030_ (.A1(_0362_),
    .A2(net28),
    .B(_0518_),
    .ZN(_0095_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1031_ (.A1(\sunrise_digital_top_i.rw_regs[38] ),
    .A2(net28),
    .ZN(_0519_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1032_ (.A1(_0365_),
    .A2(net28),
    .B(_0519_),
    .ZN(_0096_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1033_ (.A1(\sunrise_digital_top_i.rw_regs[39] ),
    .A2(net28),
    .ZN(_0520_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1034_ (.A1(_0368_),
    .A2(net28),
    .B(_0520_),
    .ZN(_0097_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1035_ (.A1(_0331_),
    .A2(_0390_),
    .Z(_0521_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1036_ (.A1(\sunrise_digital_top_i.rw_regs[40] ),
    .A2(net26),
    .ZN(_0522_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1037_ (.A1(_0344_),
    .A2(net26),
    .B(_0522_),
    .ZN(_0098_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1038_ (.A1(\sunrise_digital_top_i.rw_regs[41] ),
    .A2(net26),
    .ZN(_0523_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1039_ (.A1(_0347_),
    .A2(net27),
    .B(_0523_),
    .ZN(_0099_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1040_ (.A1(\sunrise_digital_top_i.rw_regs[42] ),
    .A2(net26),
    .ZN(_0524_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1041_ (.A1(_0351_),
    .A2(net26),
    .B(_0524_),
    .ZN(_0100_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1042_ (.A1(\sunrise_digital_top_i.rw_regs[43] ),
    .A2(net27),
    .ZN(_0525_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1043_ (.A1(_0355_),
    .A2(net27),
    .B(_0525_),
    .ZN(_0101_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1044_ (.A1(\sunrise_digital_top_i.rw_regs[44] ),
    .A2(net27),
    .ZN(_0526_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1045_ (.A1(_0359_),
    .A2(net27),
    .B(_0526_),
    .ZN(_0102_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1046_ (.A1(\sunrise_digital_top_i.rw_regs[45] ),
    .A2(net27),
    .ZN(_0527_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1047_ (.A1(_0362_),
    .A2(net26),
    .B(_0527_),
    .ZN(_0103_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1048_ (.A1(\sunrise_digital_top_i.rw_regs[46] ),
    .A2(net26),
    .ZN(_0528_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1049_ (.A1(_0365_),
    .A2(net26),
    .B(_0528_),
    .ZN(_0104_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1050_ (.A1(\sunrise_digital_top_i.rw_regs[47] ),
    .A2(net26),
    .ZN(_0529_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1051_ (.A1(_0368_),
    .A2(net26),
    .B(_0529_),
    .ZN(_0105_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1052_ (.A1(_0331_),
    .A2(_0375_),
    .Z(_0530_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1053_ (.A1(\sunrise_digital_top_i.rw_regs[24] ),
    .A2(net24),
    .ZN(_0531_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1054_ (.A1(_0344_),
    .A2(net24),
    .B(_0531_),
    .ZN(_0106_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1055_ (.A1(_0348_),
    .A2(net24),
    .ZN(_0532_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1056_ (.A1(_0198_),
    .A2(net25),
    .B(_0532_),
    .ZN(_0107_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1057_ (.A1(\sunrise_digital_top_i.rw_regs[26] ),
    .A2(net25),
    .ZN(_0533_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1058_ (.A1(_0351_),
    .A2(net24),
    .B(_0533_),
    .ZN(_0108_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1059_ (.A1(_0356_),
    .A2(net25),
    .ZN(_0534_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1060_ (.A1(_0202_),
    .A2(net25),
    .B(_0534_),
    .ZN(_0109_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1061_ (.A1(\sunrise_digital_top_i.rw_regs[28] ),
    .A2(net25),
    .ZN(_0535_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1062_ (.A1(_0359_),
    .A2(net25),
    .B(_0535_),
    .ZN(_0110_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1063_ (.A1(\sunrise_digital_top_i.rw_regs[29] ),
    .A2(net24),
    .ZN(_0536_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1064_ (.A1(_0362_),
    .A2(net24),
    .B(_0536_),
    .ZN(_0111_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1065_ (.A1(\sunrise_digital_top_i.rw_regs[30] ),
    .A2(net24),
    .ZN(_0537_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1066_ (.A1(_0365_),
    .A2(net24),
    .B(_0537_),
    .ZN(_0112_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1067_ (.A1(\sunrise_digital_top_i.rw_regs[31] ),
    .A2(net24),
    .ZN(_0538_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1068_ (.A1(_0368_),
    .A2(net24),
    .B(_0538_),
    .ZN(_0113_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1069_ (.A1(_0331_),
    .A2(_0386_),
    .ZN(_0539_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1070_ (.A1(\sunrise_digital_top_i.rw_regs[48] ),
    .A2(net22),
    .ZN(_0540_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1071_ (.A1(_0344_),
    .A2(net22),
    .B(_0540_),
    .ZN(_0114_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1072_ (.A1(\sunrise_digital_top_i.rw_regs[49] ),
    .A2(net23),
    .ZN(_0541_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1073_ (.A1(_0347_),
    .A2(net23),
    .B(_0541_),
    .ZN(_0115_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1074_ (.A1(\sunrise_digital_top_i.rw_regs[50] ),
    .A2(net22),
    .ZN(_0542_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1075_ (.A1(_0351_),
    .A2(net22),
    .B(_0542_),
    .ZN(_0116_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1076_ (.A1(\sunrise_digital_top_i.rw_regs[51] ),
    .A2(net23),
    .ZN(_0543_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1077_ (.A1(_0355_),
    .A2(net23),
    .B(_0543_),
    .ZN(_0117_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1078_ (.A1(\sunrise_digital_top_i.rw_regs[52] ),
    .A2(net23),
    .ZN(_0544_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1079_ (.A1(_0359_),
    .A2(net23),
    .B(_0544_),
    .ZN(_0118_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1080_ (.A1(\sunrise_digital_top_i.rw_regs[53] ),
    .A2(net22),
    .ZN(_0545_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1081_ (.A1(_0362_),
    .A2(net22),
    .B(_0545_),
    .ZN(_0119_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1082_ (.A1(\sunrise_digital_top_i.rw_regs[54] ),
    .A2(net22),
    .ZN(_0546_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1083_ (.A1(_0365_),
    .A2(net22),
    .B(_0546_),
    .ZN(_0120_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1084_ (.A1(\sunrise_digital_top_i.rw_regs[55] ),
    .A2(net22),
    .ZN(_0547_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1085_ (.A1(_0368_),
    .A2(net22),
    .B(_0547_),
    .ZN(_0121_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1086_ (.A1(_0331_),
    .A2(net93),
    .Z(_0548_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1087_ (.A1(\sunrise_digital_top_i.rw_regs[16] ),
    .A2(net20),
    .ZN(_0549_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1088_ (.A1(_0344_),
    .A2(net20),
    .B(_0549_),
    .ZN(_0122_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1089_ (.A1(\sunrise_digital_top_i.rw_regs[17] ),
    .A2(net20),
    .ZN(_0550_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1090_ (.A1(_0347_),
    .A2(net21),
    .B(_0550_),
    .ZN(_0123_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1091_ (.A1(\sunrise_digital_top_i.rw_regs[18] ),
    .A2(net20),
    .ZN(_0551_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1092_ (.A1(_0351_),
    .A2(net20),
    .B(_0551_),
    .ZN(_0124_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1093_ (.A1(\sunrise_digital_top_i.rw_regs[19] ),
    .A2(net21),
    .ZN(_0552_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1094_ (.A1(_0355_),
    .A2(net21),
    .B(_0552_),
    .ZN(_0125_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1095_ (.A1(\sunrise_digital_top_i.rw_regs[20] ),
    .A2(net21),
    .ZN(_0553_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1096_ (.A1(_0359_),
    .A2(net21),
    .B(_0553_),
    .ZN(_0126_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1097_ (.A1(\sunrise_digital_top_i.rw_regs[21] ),
    .A2(net21),
    .ZN(_0554_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1098_ (.A1(_0362_),
    .A2(net20),
    .B(_0554_),
    .ZN(_0127_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1099_ (.A1(\sunrise_digital_top_i.rw_regs[22] ),
    .A2(net20),
    .ZN(_0555_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1100_ (.A1(_0365_),
    .A2(net20),
    .B(_0555_),
    .ZN(_0128_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1101_ (.A1(\sunrise_digital_top_i.rw_regs[23] ),
    .A2(net20),
    .ZN(_0556_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1102_ (.A1(_0368_),
    .A2(net20),
    .B(_0556_),
    .ZN(_0129_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1103_ (.A1(_0331_),
    .A2(_0389_),
    .Z(_0557_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1104_ (.A1(\sunrise_digital_top_i.rw_regs[8] ),
    .A2(net18),
    .ZN(_0558_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1105_ (.A1(_0344_),
    .A2(net18),
    .B(_0558_),
    .ZN(_0130_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1106_ (.A1(\sunrise_digital_top_i.rw_regs[9] ),
    .A2(net18),
    .ZN(_0559_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1107_ (.A1(_0347_),
    .A2(net19),
    .B(_0559_),
    .ZN(_0131_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1108_ (.A1(\sunrise_digital_top_i.rw_regs[10] ),
    .A2(net18),
    .ZN(_0560_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1109_ (.A1(_0351_),
    .A2(net18),
    .B(_0560_),
    .ZN(_0132_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1110_ (.A1(\sunrise_digital_top_i.rw_regs[11] ),
    .A2(net19),
    .ZN(_0561_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1111_ (.A1(_0355_),
    .A2(net19),
    .B(_0561_),
    .ZN(_0133_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1112_ (.A1(\sunrise_digital_top_i.rw_regs[12] ),
    .A2(net19),
    .ZN(_0562_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1113_ (.A1(_0359_),
    .A2(net19),
    .B(_0562_),
    .ZN(_0134_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1114_ (.A1(\sunrise_digital_top_i.rw_regs[13] ),
    .A2(net19),
    .ZN(_0563_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1115_ (.A1(_0362_),
    .A2(net18),
    .B(_0563_),
    .ZN(_0135_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1116_ (.A1(\sunrise_digital_top_i.rw_regs[14] ),
    .A2(net18),
    .ZN(_0564_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1117_ (.A1(_0365_),
    .A2(net18),
    .B(_0564_),
    .ZN(_0136_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1118_ (.A1(\sunrise_digital_top_i.rw_regs[15] ),
    .A2(net18),
    .ZN(_0565_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1119_ (.A1(_0368_),
    .A2(net18),
    .B(_0565_),
    .ZN(_0137_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1120_ (.A1(_0331_),
    .A2(net40),
    .ZN(_0566_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1121_ (.A1(\sunrise_digital_top_i.rw_regs[0] ),
    .A2(net16),
    .ZN(_0567_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1122_ (.A1(_0344_),
    .A2(net16),
    .B(_0567_),
    .ZN(_0138_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1123_ (.A1(\sunrise_digital_top_i.rw_regs[1] ),
    .A2(net17),
    .ZN(_0568_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1124_ (.A1(_0347_),
    .A2(net17),
    .B(_0568_),
    .ZN(_0139_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1125_ (.A1(\sunrise_digital_top_i.rw_regs[2] ),
    .A2(net16),
    .ZN(_0569_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1126_ (.A1(_0351_),
    .A2(net16),
    .B(_0569_),
    .ZN(_0140_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1127_ (.A1(\sunrise_digital_top_i.rw_regs[3] ),
    .A2(net17),
    .ZN(_0570_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1128_ (.A1(_0355_),
    .A2(net17),
    .B(_0570_),
    .ZN(_0141_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1129_ (.A1(\sunrise_digital_top_i.rw_regs[4] ),
    .A2(net17),
    .ZN(_0571_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1130_ (.A1(_0359_),
    .A2(net17),
    .B(_0571_),
    .ZN(_0142_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1131_ (.A1(\sunrise_digital_top_i.rw_regs[5] ),
    .A2(net16),
    .ZN(_0572_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1132_ (.A1(_0362_),
    .A2(net16),
    .B(_0572_),
    .ZN(_0143_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1133_ (.A1(\sunrise_digital_top_i.rw_regs[6] ),
    .A2(net16),
    .ZN(_0573_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1134_ (.A1(_0365_),
    .A2(net16),
    .B(_0573_),
    .ZN(_0144_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1135_ (.A1(\sunrise_digital_top_i.rw_regs[7] ),
    .A2(net16),
    .ZN(_0574_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1136_ (.A1(_0368_),
    .A2(net16),
    .B(_0574_),
    .ZN(_0145_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1137_ (.A1(_0247_),
    .A2(_0259_),
    .A3(_0270_),
    .ZN(_0575_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1138_ (.A1(net30),
    .A2(_0575_),
    .ZN(_0576_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1139_ (.A1(_0260_),
    .A2(_0271_),
    .B1(net30),
    .B2(_0218_),
    .C(_0576_),
    .ZN(_0577_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1140_ (.A1(net30),
    .A2(_0577_),
    .ZN(_0578_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1141_ (.A1(net30),
    .A2(_0577_),
    .B(_0028_),
    .ZN(_0579_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1142_ (.A1(_0028_),
    .A2(net11),
    .B(_0579_),
    .ZN(_0146_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1143_ (.A1(_0028_),
    .A2(net11),
    .B(_0029_),
    .ZN(_0580_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1144_ (.A1(_0028_),
    .A2(_0029_),
    .ZN(_0581_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1145_ (.A1(net30),
    .A2(_0581_),
    .ZN(_0582_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1146_ (.A1(net11),
    .A2(_0582_),
    .B(_0580_),
    .ZN(_0147_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1147_ (.A1(_0028_),
    .A2(_0029_),
    .A3(_0030_),
    .ZN(_0583_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1148_ (.A1(_0209_),
    .A2(_0581_),
    .ZN(_0584_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1149_ (.A1(net30),
    .A2(_0583_),
    .A3(_0584_),
    .Z(_0585_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1150_ (.I0(_0030_),
    .I1(_0585_),
    .S(net11),
    .Z(_0148_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1151_ (.A1(_0591_),
    .A2(_0583_),
    .Z(_0586_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1152_ (.A1(_0183_),
    .A2(_0577_),
    .B1(_0578_),
    .B2(_0586_),
    .ZN(_0149_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1153_ (.A1(net68),
    .A2(\sunrise_digital_top_i.sync_input_spi_cs_n.data_sync[1] ),
    .ZN(_0587_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1154_ (.A1(net71),
    .A2(_0175_),
    .B(_0587_),
    .ZN(_0150_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1155_ (.I0(\sunrise_digital_top_i.sync_input_spi_mosi.data_sync[1] ),
    .I1(net10),
    .S(net68),
    .Z(_0151_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1156_ (.A1(net68),
    .A2(\sunrise_digital_top_i.sync_input_prot_sel.data_sync[1] ),
    .ZN(_0588_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1157_ (.A1(net68),
    .A2(_0191_),
    .B(_0588_),
    .ZN(_0152_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1158_ (.I0(\sunrise_digital_top_i.sync_input_spi_clk.data_sync[1] ),
    .I1(net9),
    .S(net68),
    .Z(_0153_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1159_ (.I0(\sunrise_digital_top_i.cpol_sync ),
    .I1(\sunrise_digital_top_i.sync_input_spi_cpol.data_sync[1] ),
    .S(net70),
    .Z(_0154_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1160_ (.A1(net68),
    .A2(\sunrise_digital_top_i.sync_input_spi_cs_n.data_sync[1] ),
    .ZN(_0589_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1161_ (.A1(net68),
    .A2(uio_oe[3]),
    .B(_0589_),
    .ZN(_0155_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1162_ (.A1(net71),
    .A2(\sunrise_digital_top_i.sync_input_spi_clk.data_sync[1] ),
    .ZN(_0590_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1163_ (.A1(net71),
    .A2(_0194_),
    .B(_0590_),
    .ZN(_0156_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1164_ (.I0(\sunrise_digital_top_i.sync_input_spi_cpha.data_sync[1] ),
    .I1(net4),
    .S(net70),
    .Z(_0157_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1165_ (.I0(\sunrise_digital_top_i.cpha_sync ),
    .I1(\sunrise_digital_top_i.sync_input_spi_cpha.data_sync[1] ),
    .S(net70),
    .Z(_0158_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1166_ (.I0(\sunrise_digital_top_i.sync_input_spi_cpol.data_sync[1] ),
    .I1(net3),
    .S(net70),
    .Z(_0159_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1167_ (.I0(\sunrise_digital_top_i.sync_input_prot_sel.data_sync[1] ),
    .I1(net5),
    .S(net71),
    .Z(_0160_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _1168_ (.D(_0011_),
    .SETN(net65),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1169_ (.D(_0012_),
    .RN(net64),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1170_ (.D(_0013_),
    .RN(net64),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1171_ (.D(_0014_),
    .RN(net64),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1172_ (.D(_0015_),
    .RN(net65),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.state[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1173_ (.D(_0031_),
    .RN(net64),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_spi_clk.data_dly ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1174_ (.D(_0000_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0161_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1175_ (.D(_0001_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0162_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1176_ (.D(_0002_),
    .RN(net51),
    .CLK(clknet_4_5_0_clk),
    .Q(_0163_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1177_ (.D(_0003_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0164_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1178_ (.D(_0004_),
    .RN(net51),
    .CLK(clknet_4_5_0_clk),
    .Q(_0165_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1179_ (.D(_0005_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0166_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1180_ (.D(_0006_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0167_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1181_ (.D(_0007_),
    .RN(net52),
    .CLK(clknet_4_5_0_clk),
    .Q(_0168_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1182_ (.D(_0008_),
    .RN(net52),
    .CLK(clknet_4_5_0_clk),
    .Q(_0169_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1183_ (.D(_0032_),
    .RN(net64),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.falling_edge_detector_sof.data_dly ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1184_ (.D(_0033_),
    .RN(net60),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1185_ (.D(_0034_),
    .RN(net60),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1186_ (.D(_0035_),
    .RN(net60),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1187_ (.D(_0036_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1188_ (.D(_0037_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1189_ (.D(_0038_),
    .RN(net63),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1190_ (.D(_0039_),
    .RN(net65),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1191_ (.D(_0040_),
    .RN(net65),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1192_ (.D(_0041_),
    .RN(net60),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1193_ (.D(_0042_),
    .RN(net60),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1194_ (.D(_0043_),
    .RN(net60),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1195_ (.D(_0044_),
    .RN(net64),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1196_ (.D(_0045_),
    .RN(net64),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[17] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1197_ (.D(_0046_),
    .RN(net65),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.mux_addr_i.a[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1198_ (.D(_0047_),
    .RN(net65),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1199_ (.D(_0048_),
    .RN(net65),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1200_ (.D(_0049_),
    .RN(net65),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1201_ (.D(_0050_),
    .RN(net65),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.buffer_counter[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1202_ (.D(_0051_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[56] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1203_ (.D(_0052_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[57] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1204_ (.D(_0053_),
    .RN(net53),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[58] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1205_ (.D(_0054_),
    .RN(net63),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[59] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1206_ (.D(_0055_),
    .RN(net63),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[60] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1207_ (.D(_0056_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[61] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1208_ (.D(_0057_),
    .RN(net54),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[62] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1209_ (.D(_0058_),
    .RN(net49),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[63] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1210_ (.D(_0059_),
    .RN(net60),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1211_ (.D(_0060_),
    .RN(net60),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1212_ (.D(_0061_),
    .RN(net62),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1213_ (.D(_0062_),
    .RN(net62),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1214_ (.D(_0063_),
    .RN(net62),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1215_ (.D(_0064_),
    .RN(net62),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1216_ (.D(_0065_),
    .RN(net55),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.tx_buffer[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1217_ (.D(_0066_),
    .RN(net55),
    .CLK(clknet_4_7_0_clk),
    .Q(spi_miso),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1218_ (.D(_0067_),
    .RN(net61),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1219_ (.D(_0068_),
    .RN(net64),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1220_ (.D(_0069_),
    .RN(net64),
    .CLK(clknet_4_14_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1221_ (.D(_0070_),
    .RN(net64),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1222_ (.D(_0071_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1223_ (.D(_0072_),
    .RN(net67),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1224_ (.D(_0073_),
    .RN(net67),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1225_ (.D(_0074_),
    .RN(net65),
    .CLK(clknet_4_11_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.spi_peripheral_i.rx_buffer[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1226_ (.D(_0009_),
    .CLK(clknet_4_5_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1227_ (.D(_0010_),
    .CLK(clknet_4_5_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.last_event[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1228_ (.D(_0017_),
    .RN(net52),
    .CLK(clknet_4_5_0_clk),
    .Q(_0024_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 _1229_ (.D(_0018_),
    .RN(net52),
    .CLK(clknet_4_5_0_clk),
    .Q(_0025_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1230_ (.D(_0019_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0026_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1231_ (.D(_0020_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(_0027_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1232_ (.D(_0075_),
    .RN(net55),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1233_ (.D(_0076_),
    .RN(net55),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1234_ (.D(_0077_),
    .RN(net62),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1235_ (.D(_0078_),
    .RN(net62),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1236_ (.D(_0079_),
    .RN(net55),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1237_ (.D(_0080_),
    .RN(net55),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1238_ (.D(_0081_),
    .RN(net56),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1239_ (.D(_0082_),
    .RN(net52),
    .CLK(clknet_4_5_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.pull_sda ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1240_ (.D(_0083_),
    .RN(net55),
    .CLK(clknet_4_6_0_clk),
    .Q(_0016_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1241_ (.D(_0084_),
    .RN(net55),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1242_ (.D(_0085_),
    .RN(net56),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1243_ (.D(_0086_),
    .RN(net56),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1244_ (.D(_0087_),
    .RN(net62),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_addr[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1245_ (.D(_0021_),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_start ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1246_ (.D(_0023_),
    .RN(net51),
    .CLK(clknet_4_4_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.we ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1247_ (.D(_0022_),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.bus_stop ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1248_ (.D(_0088_),
    .RN(net61),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.spi_mosi_sync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1249_ (.D(net6),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1250_ (.D(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[0] ),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1251_ (.D(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[1] ),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1252_ (.D(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[2] ),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.sda_d[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1253_ (.D(_0089_),
    .RN(net55),
    .CLK(clknet_4_6_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.dbyte[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1254_ (.D(net7),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1255_ (.D(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[0] ),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1256_ (.D(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[1] ),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1257_ (.D(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[2] ),
    .CLK(clknet_4_7_0_clk),
    .Q(\sunrise_digital_top_i.top_wrapper_i.i2c_peripheral_i.scl_d[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1258_ (.D(_0090_),
    .RN(net54),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[32] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1259_ (.D(_0091_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[33] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1260_ (.D(_0092_),
    .RN(net53),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[34] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1261_ (.D(_0093_),
    .RN(net59),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[35] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1262_ (.D(_0094_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[36] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1263_ (.D(_0095_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[37] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1264_ (.D(_0096_),
    .RN(net54),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[38] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1265_ (.D(_0097_),
    .RN(net54),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[39] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1266_ (.D(_0098_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[40] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1267_ (.D(_0099_),
    .RN(net58),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[41] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1268_ (.D(_0100_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[42] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1269_ (.D(_0101_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[43] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1270_ (.D(_0102_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[44] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1271_ (.D(_0103_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[45] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1272_ (.D(_0104_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[46] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1273_ (.D(_0105_),
    .RN(net49),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[47] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1274_ (.D(_0106_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[24] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1275_ (.D(_0107_),
    .RN(net59),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[25] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1276_ (.D(_0108_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[26] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1277_ (.D(_0109_),
    .RN(net59),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[27] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1278_ (.D(_0110_),
    .RN(net59),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[28] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1279_ (.D(_0111_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[29] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1280_ (.D(_0112_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[30] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1281_ (.D(_0113_),
    .RN(net49),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[31] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1282_ (.D(_0114_),
    .RN(net54),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[48] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1283_ (.D(_0115_),
    .RN(net58),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[49] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1284_ (.D(_0116_),
    .RN(net53),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[50] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1285_ (.D(_0117_),
    .RN(net59),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[51] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1286_ (.D(_0118_),
    .RN(net59),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[52] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1287_ (.D(_0119_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[53] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1288_ (.D(_0120_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[54] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1289_ (.D(_0121_),
    .RN(net54),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[55] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1290_ (.D(_0122_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[16] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1291_ (.D(_0123_),
    .RN(net63),
    .CLK(clknet_4_10_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[17] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1292_ (.D(_0124_),
    .RN(net53),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[18] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1293_ (.D(_0125_),
    .RN(net59),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[19] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1294_ (.D(_0126_),
    .RN(net59),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[20] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1295_ (.D(_0127_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[21] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1296_ (.D(_0128_),
    .RN(net49),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[22] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1297_ (.D(_0129_),
    .RN(net50),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[23] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1298_ (.D(_0130_),
    .RN(net54),
    .CLK(clknet_4_0_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1299_ (.D(_0131_),
    .RN(net58),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1300_ (.D(_0132_),
    .RN(net56),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1301_ (.D(_0133_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1302_ (.D(_0134_),
    .RN(net67),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1303_ (.D(_0135_),
    .RN(net58),
    .CLK(clknet_4_8_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1304_ (.D(_0136_),
    .RN(net54),
    .CLK(clknet_4_2_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1305_ (.D(_0137_),
    .RN(net50),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1306_ (.D(_0138_),
    .RN(net54),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1307_ (.D(_0139_),
    .RN(net60),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1308_ (.D(_0140_),
    .RN(net56),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1309_ (.D(_0141_),
    .RN(net67),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1310_ (.D(_0142_),
    .RN(net59),
    .CLK(clknet_4_9_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1311_ (.D(_0143_),
    .RN(net56),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1312_ (.D(_0144_),
    .RN(net55),
    .CLK(clknet_4_3_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1313_ (.D(_0145_),
    .RN(net54),
    .CLK(clknet_4_1_0_clk),
    .Q(\sunrise_digital_top_i.rw_regs[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1314_ (.D(_0146_),
    .RN(net50),
    .CLK(clknet_4_1_0_clk),
    .Q(_0028_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1315_ (.D(_0147_),
    .RN(net50),
    .CLK(clknet_4_1_0_clk),
    .Q(_0029_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1316_ (.D(_0148_),
    .RN(net50),
    .CLK(clknet_4_1_0_clk),
    .Q(_0030_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1317_ (.D(_0149_),
    .RN(net57),
    .CLK(clknet_4_4_0_clk),
    .Q(_0591_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1318_ (.D(_0150_),
    .RN(net61),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.spi_cs_n_sync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1319_ (.D(_0151_),
    .RN(net62),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.sync_input_spi_mosi.data_sync[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _1320_ (.D(_0152_),
    .RN(net60),
    .CLK(clknet_4_12_0_clk),
    .Q(\sunrise_digital_top_i.protrocol_sel_sync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1321_ (.D(_0153_),
    .RN(net61),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.sync_input_spi_clk.data_sync[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1322_ (.D(_0154_),
    .RN(net66),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.cpol_sync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1323_ (.D(_0155_),
    .RN(net61),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.sync_input_spi_cs_n.data_sync[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1324_ (.D(_0156_),
    .RN(net66),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.spi_clk_sync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1325_ (.D(_0157_),
    .RN(net66),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.sync_input_spi_cpha.data_sync[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1326_ (.D(_0158_),
    .RN(net66),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.cpha_sync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1327_ (.D(_0159_),
    .RN(net66),
    .CLK(clknet_4_15_0_clk),
    .Q(\sunrise_digital_top_i.sync_input_spi_cpol.data_sync[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _1328_ (.D(_0160_),
    .RN(net61),
    .CLK(clknet_4_13_0_clk),
    .Q(\sunrise_digital_top_i.sync_input_prot_sel.data_sync[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_73 (.ZN(net73),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_74 (.ZN(net74),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_75 (.ZN(net75),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_76 (.ZN(net76),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_77 (.ZN(net77),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_78 (.ZN(net78),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_79 (.ZN(net79),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_80 (.ZN(net80),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_81 (.ZN(net81),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_82 (.ZN(net82),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_83 (.ZN(net83),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_84 (.ZN(net84),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_85 (.ZN(net85),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_86 (.ZN(net86),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_87 (.ZN(net87),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_88 (.ZN(net88),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_89 (.ZN(net89),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_90 (.ZN(net90),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_91 (.ZN(net91),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_92 (.ZN(net92),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1350_ (.I(i2c_sda_oe),
    .Z(uio_oe[1]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _1351_ (.I(spi_miso),
    .Z(uio_out[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_39 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_40 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_41 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_42 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_43 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_44 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_45 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_46 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_47 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_48 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_49 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_50 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_51 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_52 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_53 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_54 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_55 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_56 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_57 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_58 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_59 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_60 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_61 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_62 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_63 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_64 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_65 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_66 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_67 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_68 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_69 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_70 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_71 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_72 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_73 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_74 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_75 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_76 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_77 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_78 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_79 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_80 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_81 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_82 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_83 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_84 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_85 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_86 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_87 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_88 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_89 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_95 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_96 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_97 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_98 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_99 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_103 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_109 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_110 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_111 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_113 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_114 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_115 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_116 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_117 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_118 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_119 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_120 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_121 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_122 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_123 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_124 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_125 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_126 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_127 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_128 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_129 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_130 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_131 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_132 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_133 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_134 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_135 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_136 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_137 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_138 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_139 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_140 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_141 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_142 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_143 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_144 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_145 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_146 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_147 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_148 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_149 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_150 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_151 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_152 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_153 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_154 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_155 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_156 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_157 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_158 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_159 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_160 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_161 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_162 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_163 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_164 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_165 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_166 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_167 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_168 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_169 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_170 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_171 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_172 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_173 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_174 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_175 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_176 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_177 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_178 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_179 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_180 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_181 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_182 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_183 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_184 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_185 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_186 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_187 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_188 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_189 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_190 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_191 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_192 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_193 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_194 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_195 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_196 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_197 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_198 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_199 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_200 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_201 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_202 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_203 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_204 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_205 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_206 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_207 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_208 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_209 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_210 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_211 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_212 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_213 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_214 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_215 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_216 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_217 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_218 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_219 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_220 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_221 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_222 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_223 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_224 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_225 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_226 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_227 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_228 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_229 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_230 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_231 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_232 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_233 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_234 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_235 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_236 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_237 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_238 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_239 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_240 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_241 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_242 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_243 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_244 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_245 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_246 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_247 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_248 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_249 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_250 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_251 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_252 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_253 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_254 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_255 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_256 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_257 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_258 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_259 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_260 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_261 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_262 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_263 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_264 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_265 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_266 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_267 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_268 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_269 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_270 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_271 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_272 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_273 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_274 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_275 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_276 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_277 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_278 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_279 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_280 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_281 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_282 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_283 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_284 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_285 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_286 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_287 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_288 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_289 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_290 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_291 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_292 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_293 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_294 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_295 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_296 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_297 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_298 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_299 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_300 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_301 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_302 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_303 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_304 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_305 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_306 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_307 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_308 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_309 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_310 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_311 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_312 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_313 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_314 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_315 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_316 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_317 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_318 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_319 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_320 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_321 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_322 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_323 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_324 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_325 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_326 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_327 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_328 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_329 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_330 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_331 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_332 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_333 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_334 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_335 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_336 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_337 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_338 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_339 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_340 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_341 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_342 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_343 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_344 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_345 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_346 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_347 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_348 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_349 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_350 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_351 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_352 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_353 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_354 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_355 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_356 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_357 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_358 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_359 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_360 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_361 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_362 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_363 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_364 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_365 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_366 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_367 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_368 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_369 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_370 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_371 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_372 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_373 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_374 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_375 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_376 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_377 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_378 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_379 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_380 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_381 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_382 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_383 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_384 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_385 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_386 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_387 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_388 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_389 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_390 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_391 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_392 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_393 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_394 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_395 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_396 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_397 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_398 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_399 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_400 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_401 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_402 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_403 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_404 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_405 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_406 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_407 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_409 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_410 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_411 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_412 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_413 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_414 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_416 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_417 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_418 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_419 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_420 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_421 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_422 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_423 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_424 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_425 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(ena),
    .Z(net1),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(rst_n),
    .Z(net2),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(ui_in[0]),
    .Z(net3),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(ui_in[1]),
    .Z(net4),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(ui_in[7]),
    .Z(net5),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(uio_in[1]),
    .Z(net6),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(uio_in[2]),
    .Z(net7),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(uio_in[4]),
    .Z(net8),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(uio_in[5]),
    .Z(net9),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(uio_in[6]),
    .Z(net10),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 max_cap11 (.I(_0577_),
    .Z(net11),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout12 (.I(_0469_),
    .Z(net12),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 max_cap13 (.I(_0451_),
    .Z(net13),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 max_cap14 (.I(_0443_),
    .Z(net14),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout15 (.I(_0282_),
    .Z(net15),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout16 (.I(_0566_),
    .Z(net16),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout17 (.I(_0566_),
    .Z(net17),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout18 (.I(_0557_),
    .Z(net18),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout19 (.I(_0557_),
    .Z(net19),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout20 (.I(_0548_),
    .Z(net20),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout21 (.I(_0548_),
    .Z(net21),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout22 (.I(_0539_),
    .Z(net22),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout23 (.I(_0539_),
    .Z(net23),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout24 (.I(_0530_),
    .Z(net24),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout25 (.I(_0530_),
    .Z(net25),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout26 (.I(_0521_),
    .Z(net26),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout27 (.I(_0521_),
    .Z(net27),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout28 (.I(_0512_),
    .Z(net28),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout29 (.I(_0512_),
    .Z(net29),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout30 (.I(_0471_),
    .Z(net30),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 wire32 (.I(_0428_),
    .Z(net32),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 wire33 (.I(_0420_),
    .Z(net33),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 wire34 (.I(_0400_),
    .Z(net34),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout35 (.I(_0342_),
    .Z(net35),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout36 (.I(_0342_),
    .Z(net36),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout37 (.I(_0322_),
    .Z(net37),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 wire38 (.I(_0421_),
    .Z(net38),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout39 (.I(_0383_),
    .Z(net39),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout40 (.I(_0383_),
    .Z(net40),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout41 (.I(_0377_),
    .Z(net41),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 max_cap42 (.I(_0243_),
    .Z(net42),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout43 (.I(_0215_),
    .Z(net43),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout44 (.I(_0340_),
    .Z(net44),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout45 (.I(_0335_),
    .Z(net45),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout46 (.I(net48),
    .Z(net46),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout47 (.I(net48),
    .Z(net47),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 fanout48 (.I(\sunrise_digital_top_i.protrocol_sel_sync ),
    .Z(net48),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout49 (.I(net50),
    .Z(net49),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout50 (.I(net57),
    .Z(net50),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout51 (.I(net57),
    .Z(net51),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout52 (.I(net57),
    .Z(net52),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout53 (.I(net56),
    .Z(net53),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout54 (.I(net56),
    .Z(net54),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout55 (.I(net56),
    .Z(net55),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout56 (.I(net57),
    .Z(net56),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout57 (.I(net2),
    .Z(net57),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout58 (.I(net59),
    .Z(net58),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout59 (.I(net67),
    .Z(net59),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout60 (.I(net62),
    .Z(net60),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout61 (.I(net62),
    .Z(net61),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout62 (.I(net67),
    .Z(net62),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout63 (.I(net67),
    .Z(net63),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout64 (.I(net66),
    .Z(net64),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout65 (.I(net66),
    .Z(net65),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout66 (.I(net67),
    .Z(net66),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout67 (.I(net2),
    .Z(net67),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout68 (.I(net71),
    .Z(net68),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 fanout69 (.I(net71),
    .Z(net69),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout70 (.I(net71),
    .Z(net70),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout71 (.I(net1),
    .Z(net71),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__tiel tt_um_calonso88_spi_i2c_reg_bank_72 (.ZN(net72),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload0 (.I(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload1 (.I(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkload2 (.I(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload3 (.I(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload4 (.I(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload5 (.I(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload6 (.I(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 clkload7 (.I(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload8 (.I(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload9 (.I(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload10 (.I(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload11 (.I(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload12 (.I(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload13 (.I(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 clone1 (.A1(_0339_),
    .A2(net95),
    .Z(net93),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer2 (.I(_0385_),
    .Z(net94),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer3 (.I(net94),
    .Z(net95),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer4 (.I(_0385_),
    .Z(net96),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer5 (.I(net48),
    .Z(net97),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer6 (.I(net97),
    .Z(net98),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_316 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_326 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_334 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_596 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_166 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_168 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_218 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_230 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_238 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_287 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_299 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_334 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_456 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_294 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_371 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_403 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_497 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_200 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_297 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_366 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_414 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_435 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_471 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_487 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_256 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_264 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_328 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_336 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_401 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_433 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_441 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_443 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_188 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_196 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_218 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_250 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_266 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_334 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_373 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_377 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_441 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_167 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_229 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_281 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_289 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_367 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_406 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_471 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_509 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_217 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_270 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_363 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_371 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_375 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_234 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_258 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_299 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_335 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_391 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_437 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_511 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_519 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_176 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_214 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_237 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_253 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_315 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_414 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_438 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_442 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_232 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_236 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_332 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_365 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_367 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_516 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_217 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_299 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_305 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_374 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_466 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_487 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_187 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_373 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_445 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_196 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_198 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_218 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_310 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_328 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_330 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_442 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_502 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_537 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_553 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_214 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_229 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_463 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_471 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_475 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_574 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_166 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_218 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_250 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_266 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_284 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_386 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_396 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_181 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_237 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_305 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_351 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_368 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_583 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_201 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_551 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_596 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_115 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_184 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_200 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_210 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_261 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_265 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_355 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_392 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_394 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_415 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_440 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_472 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_503 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_519 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_535 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_573 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_589 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_187 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_222 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_270 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_310 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_438 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_526 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_596 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_123 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_213 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_272 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_305 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_472 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_476 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_560 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_88 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_92 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_166 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_170 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_200 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_228 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_236 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_345 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_437 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_441 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_443 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_507 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_515 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_551 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_126 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_161 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_169 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_232 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_258 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_262 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_351 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_367 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_403 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_445 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_499 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_515 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_561 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_569 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_88 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_135 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_272 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_310 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_327 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_467 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_483 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_487 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_504 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_506 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_541 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_550 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_566 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_77 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_81 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_83 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_88 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_120 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_144 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_305 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_378 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_403 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_411 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_449 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_537 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_545 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_549 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_133 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_297 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_299 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_332 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_401 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_477 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_550 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_554 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_61 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_65 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_102 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_391 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_540 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_560 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_589 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_88 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_270 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_407 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_472 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_515 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_553 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_61 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_99 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_290 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_344 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_350 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_364 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_445 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_479 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_516 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_518 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_246 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_316 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_369 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_373 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_409 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_438 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_477 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_501 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_509 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_599 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_603 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_85 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_228 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_351 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_359 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_363 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_433 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_437 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_514 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_566 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_575 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_80 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_246 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_248 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_327 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_61 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_65 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_112 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_123 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_190 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_287 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_297 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_357 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_363 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_459 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_491 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_501 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_509 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_578 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_88 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_92 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_94 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_129 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_170 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_183 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_237 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_288 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_364 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_375 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_426 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_480 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_484 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_507 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_120 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_144 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_159 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_168 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_211 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_283 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_287 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_340 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_380 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_400 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_435 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_443 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_471 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_475 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_531 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_585 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_120 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_245 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_305 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_335 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_390 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_392 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_458 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_466 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_468 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_548 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_577 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_601 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_115 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_165 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_200 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_210 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_214 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_319 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_466 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_516 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_162 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_362 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_434 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_541 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_600 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_604 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_36 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_52 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_57 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_65 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_74 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_78 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_83 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_91 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_96 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_100 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_112 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_130 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_134 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_161 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_169 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_176 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_180 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_182 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_187 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_200 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_214 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_237 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_252 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_265 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_335 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_350 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_372 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_394 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_475 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_539 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_571 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 assign uio_oe[0] = net72;
 assign uio_oe[2] = net73;
 assign uio_oe[4] = net74;
 assign uio_oe[5] = net75;
 assign uio_oe[6] = net76;
 assign uio_oe[7] = net77;
 assign uio_out[0] = net78;
 assign uio_out[1] = net79;
 assign uio_out[2] = net80;
 assign uio_out[4] = net81;
 assign uio_out[5] = net82;
 assign uio_out[6] = net83;
 assign uio_out[7] = net84;
 assign uo_out[0] = net85;
 assign uo_out[1] = net86;
 assign uo_out[2] = net87;
 assign uo_out[3] = net88;
 assign uo_out[4] = net89;
 assign uo_out[5] = net90;
 assign uo_out[6] = net91;
 assign uo_out[7] = net92;
endmodule

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_MichaelBell_tinyQV
  CLASS BLOCK ;
  FOREIGN tt_um_MichaelBell_tinyQV ;
  ORIGIN 0.000 0.000 ;
  SIZE 1075.760 BY 736.960 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.780 3.620 177.380 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.380 3.620 330.980 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 482.980 3.620 484.580 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.580 3.620 638.180 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.180 3.620 791.780 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.780 3.620 945.380 733.340 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.480 3.620 174.080 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.080 3.620 327.680 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 479.680 3.620 481.280 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 633.280 3.620 634.880 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 786.880 3.620 788.480 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 940.480 3.620 942.080 733.340 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 312.890 735.960 313.190 736.960 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 320.170 735.960 320.470 736.960 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 305.610 735.960 305.910 736.960 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    PORT
      LAYER Metal4 ;
        RECT 298.330 735.960 298.630 736.960 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 291.050 735.960 291.350 736.960 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 283.770 735.960 284.070 736.960 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 276.490 735.960 276.790 736.960 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 269.210 735.960 269.510 736.960 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 261.930 735.960 262.230 736.960 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 254.650 735.960 254.950 736.960 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 247.370 735.960 247.670 736.960 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 240.090 735.960 240.390 736.960 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 232.810 735.960 233.110 736.960 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 225.530 735.960 225.830 736.960 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 218.250 735.960 218.550 736.960 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 210.970 735.960 211.270 736.960 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    PORT
      LAYER Metal4 ;
        RECT 203.690 735.960 203.990 736.960 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 196.410 735.960 196.710 736.960 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 189.130 735.960 189.430 736.960 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 65.370 735.960 65.670 736.960 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.879200 ;
    PORT
      LAYER Metal4 ;
        RECT 58.090 735.960 58.390 736.960 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 50.810 735.960 51.110 736.960 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 43.530 735.960 43.830 736.960 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 36.250 735.960 36.550 736.960 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 3.879200 ;
    PORT
      LAYER Metal4 ;
        RECT 28.970 735.960 29.270 736.960 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 21.690 735.960 21.990 736.960 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 14.410 735.960 14.710 736.960 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 123.610 735.960 123.910 736.960 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.879200 ;
    PORT
      LAYER Metal4 ;
        RECT 116.330 735.960 116.630 736.960 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 109.050 735.960 109.350 736.960 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.365600 ;
    PORT
      LAYER Metal4 ;
        RECT 101.770 735.960 102.070 736.960 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.389000 ;
    PORT
      LAYER Metal4 ;
        RECT 94.490 735.960 94.790 736.960 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256000 ;
    PORT
      LAYER Metal4 ;
        RECT 87.210 735.960 87.510 736.960 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 79.930 735.960 80.230 736.960 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.389000 ;
    PORT
      LAYER Metal4 ;
        RECT 72.650 735.960 72.950 736.960 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.028900 ;
    PORT
      LAYER Metal4 ;
        RECT 181.850 735.960 182.150 736.960 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 174.570 735.960 174.870 736.960 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 167.290 735.960 167.590 736.960 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.304600 ;
    PORT
      LAYER Metal4 ;
        RECT 160.010 735.960 160.310 736.960 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 152.730 735.960 153.030 736.960 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 145.450 735.960 145.750 736.960 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 138.170 735.960 138.470 736.960 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 130.890 735.960 131.190 736.960 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 3.490 1073.390 733.470 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 1072.960 733.340 ;
      LAYER Metal2 ;
        RECT 1.820 0.650 1072.260 734.630 ;
      LAYER Metal3 ;
        RECT 1.770 0.700 1072.310 734.580 ;
      LAYER Metal4 ;
        RECT 8.540 735.660 14.110 735.960 ;
        RECT 15.010 735.660 21.390 735.960 ;
        RECT 22.290 735.660 28.670 735.960 ;
        RECT 29.570 735.660 35.950 735.960 ;
        RECT 36.850 735.660 43.230 735.960 ;
        RECT 44.130 735.660 50.510 735.960 ;
        RECT 51.410 735.660 57.790 735.960 ;
        RECT 58.690 735.660 65.070 735.960 ;
        RECT 65.970 735.660 72.350 735.960 ;
        RECT 73.250 735.660 79.630 735.960 ;
        RECT 80.530 735.660 86.910 735.960 ;
        RECT 87.810 735.660 94.190 735.960 ;
        RECT 95.090 735.660 101.470 735.960 ;
        RECT 102.370 735.660 108.750 735.960 ;
        RECT 109.650 735.660 116.030 735.960 ;
        RECT 116.930 735.660 123.310 735.960 ;
        RECT 124.210 735.660 130.590 735.960 ;
        RECT 131.490 735.660 137.870 735.960 ;
        RECT 138.770 735.660 145.150 735.960 ;
        RECT 146.050 735.660 152.430 735.960 ;
        RECT 153.330 735.660 159.710 735.960 ;
        RECT 160.610 735.660 166.990 735.960 ;
        RECT 167.890 735.660 174.270 735.960 ;
        RECT 175.170 735.660 181.550 735.960 ;
        RECT 182.450 735.660 188.830 735.960 ;
        RECT 189.730 735.660 196.110 735.960 ;
        RECT 197.010 735.660 203.390 735.960 ;
        RECT 204.290 735.660 210.670 735.960 ;
        RECT 211.570 735.660 217.950 735.960 ;
        RECT 218.850 735.660 225.230 735.960 ;
        RECT 226.130 735.660 232.510 735.960 ;
        RECT 233.410 735.660 239.790 735.960 ;
        RECT 240.690 735.660 247.070 735.960 ;
        RECT 247.970 735.660 254.350 735.960 ;
        RECT 255.250 735.660 261.630 735.960 ;
        RECT 262.530 735.660 268.910 735.960 ;
        RECT 269.810 735.660 276.190 735.960 ;
        RECT 277.090 735.660 283.470 735.960 ;
        RECT 284.370 735.660 290.750 735.960 ;
        RECT 291.650 735.660 298.030 735.960 ;
        RECT 298.930 735.660 305.310 735.960 ;
        RECT 306.210 735.660 312.590 735.960 ;
        RECT 313.490 735.660 319.870 735.960 ;
        RECT 320.770 735.660 1068.340 735.960 ;
        RECT 8.540 733.640 1068.340 735.660 ;
        RECT 8.540 3.320 18.580 733.640 ;
        RECT 20.780 3.320 21.880 733.640 ;
        RECT 24.080 3.320 172.180 733.640 ;
        RECT 174.380 3.320 175.480 733.640 ;
        RECT 177.680 3.320 325.780 733.640 ;
        RECT 327.980 3.320 329.080 733.640 ;
        RECT 331.280 3.320 479.380 733.640 ;
        RECT 481.580 3.320 482.680 733.640 ;
        RECT 484.880 3.320 632.980 733.640 ;
        RECT 635.180 3.320 636.280 733.640 ;
        RECT 638.480 3.320 786.580 733.640 ;
        RECT 788.780 3.320 789.880 733.640 ;
        RECT 792.080 3.320 940.180 733.640 ;
        RECT 942.380 3.320 943.480 733.640 ;
        RECT 945.680 3.320 1068.340 733.640 ;
        RECT 8.540 1.210 1068.340 3.320 ;
  END
END tt_um_MichaelBell_tinyQV
END LIBRARY

